/*
 * Author: neidong_fu
 * Time  : 2020/03/04
 * function: caculate sqrt(mantissa)
*/

module man_sqrt(
    // out = sqrt(in) = round(sqrt(in/(2^10)) * 2^12) 
    input [9:0] in,          // in (0,0,10)
    output reg [11:0] out   // out(0,0,12)
    );

    always@(*)begin
        case(in)
        10'd 1:out = 12'd 128;
        10'd 2:out = 12'd 181;
        10'd 3:out = 12'd 222;
        10'd 4:out = 12'd 256;
        10'd 5:out = 12'd 286;
        10'd 6:out = 12'd 314;
        10'd 7:out = 12'd 339;
        10'd 8:out = 12'd 362;
        10'd 9:out = 12'd 384;
        10'd 10:out = 12'd 405;
        10'd 11:out = 12'd 425;
        10'd 12:out = 12'd 443;
        10'd 13:out = 12'd 462;
        10'd 14:out = 12'd 479;
        10'd 15:out = 12'd 496;
        10'd 16:out = 12'd 512;
        10'd 17:out = 12'd 528;
        10'd 18:out = 12'd 543;
        10'd 19:out = 12'd 558;
        10'd 20:out = 12'd 572;
        10'd 21:out = 12'd 587;
        10'd 22:out = 12'd 600;
        10'd 23:out = 12'd 614;
        10'd 24:out = 12'd 627;
        10'd 25:out = 12'd 640;
        10'd 26:out = 12'd 653;
        10'd 27:out = 12'd 665;
        10'd 28:out = 12'd 677;
        10'd 29:out = 12'd 689;
        10'd 30:out = 12'd 701;
        10'd 31:out = 12'd 713;
        10'd 32:out = 12'd 724;
        10'd 33:out = 12'd 735;
        10'd 34:out = 12'd 746;
        10'd 35:out = 12'd 757;
        10'd 36:out = 12'd 768;
        10'd 37:out = 12'd 779;
        10'd 38:out = 12'd 789;
        10'd 39:out = 12'd 799;
        10'd 40:out = 12'd 810;
        10'd 41:out = 12'd 820;
        10'd 42:out = 12'd 830;
        10'd 43:out = 12'd 839;
        10'd 44:out = 12'd 849;
        10'd 45:out = 12'd 859;
        10'd 46:out = 12'd 868;
        10'd 47:out = 12'd 878;
        10'd 48:out = 12'd 887;
        10'd 49:out = 12'd 896;
        10'd 50:out = 12'd 905;
        10'd 51:out = 12'd 914;
        10'd 52:out = 12'd 923;
        10'd 53:out = 12'd 932;
        10'd 54:out = 12'd 941;
        10'd 55:out = 12'd 949;
        10'd 56:out = 12'd 958;
        10'd 57:out = 12'd 966;
        10'd 58:out = 12'd 975;
        10'd 59:out = 12'd 983;
        10'd 60:out = 12'd 991;
        10'd 61:out = 12'd 1000;
        10'd 62:out = 12'd 1008;
        10'd 63:out = 12'd 1016;
        10'd 64:out = 12'd 1024;
        10'd 65:out = 12'd 1032;
        10'd 66:out = 12'd 1040;
        10'd 67:out = 12'd 1048;
        10'd 68:out = 12'd 1056;
        10'd 69:out = 12'd 1063;
        10'd 70:out = 12'd 1071;
        10'd 71:out = 12'd 1079;
        10'd 72:out = 12'd 1086;
        10'd 73:out = 12'd 1094;
        10'd 74:out = 12'd 1101;
        10'd 75:out = 12'd 1109;
        10'd 76:out = 12'd 1116;
        10'd 77:out = 12'd 1123;
        10'd 78:out = 12'd 1130;
        10'd 79:out = 12'd 1138;
        10'd 80:out = 12'd 1145;
        10'd 81:out = 12'd 1152;
        10'd 82:out = 12'd 1159;
        10'd 83:out = 12'd 1166;
        10'd 84:out = 12'd 1173;
        10'd 85:out = 12'd 1180;
        10'd 86:out = 12'd 1187;
        10'd 87:out = 12'd 1194;
        10'd 88:out = 12'd 1201;
        10'd 89:out = 12'd 1208;
        10'd 90:out = 12'd 1214;
        10'd 91:out = 12'd 1221;
        10'd 92:out = 12'd 1228;
        10'd 93:out = 12'd 1234;
        10'd 94:out = 12'd 1241;
        10'd 95:out = 12'd 1248;
        10'd 96:out = 12'd 1254;
        10'd 97:out = 12'd 1261;
        10'd 98:out = 12'd 1267;
        10'd 99:out = 12'd 1274;
        10'd 100:out = 12'd 1280;
        10'd 101:out = 12'd 1286;
        10'd 102:out = 12'd 1293;
        10'd 103:out = 12'd 1299;
        10'd 104:out = 12'd 1305;
        10'd 105:out = 12'd 1312;
        10'd 106:out = 12'd 1318;
        10'd 107:out = 12'd 1324;
        10'd 108:out = 12'd 1330;
        10'd 109:out = 12'd 1336;
        10'd 110:out = 12'd 1342;
        10'd 111:out = 12'd 1349;
        10'd 112:out = 12'd 1355;
        10'd 113:out = 12'd 1361;
        10'd 114:out = 12'd 1367;
        10'd 115:out = 12'd 1373;
        10'd 116:out = 12'd 1379;
        10'd 117:out = 12'd 1385;
        10'd 118:out = 12'd 1390;
        10'd 119:out = 12'd 1396;
        10'd 120:out = 12'd 1402;
        10'd 121:out = 12'd 1408;
        10'd 122:out = 12'd 1414;
        10'd 123:out = 12'd 1420;
        10'd 124:out = 12'd 1425;
        10'd 125:out = 12'd 1431;
        10'd 126:out = 12'd 1437;
        10'd 127:out = 12'd 1442;
        10'd 128:out = 12'd 1448;
        10'd 129:out = 12'd 1454;
        10'd 130:out = 12'd 1459;
        10'd 131:out = 12'd 1465;
        10'd 132:out = 12'd 1471;
        10'd 133:out = 12'd 1476;
        10'd 134:out = 12'd 1482;
        10'd 135:out = 12'd 1487;
        10'd 136:out = 12'd 1493;
        10'd 137:out = 12'd 1498;
        10'd 138:out = 12'd 1504;
        10'd 139:out = 12'd 1509;
        10'd 140:out = 12'd 1515;
        10'd 141:out = 12'd 1520;
        10'd 142:out = 12'd 1525;
        10'd 143:out = 12'd 1531;
        10'd 144:out = 12'd 1536;
        10'd 145:out = 12'd 1541;
        10'd 146:out = 12'd 1547;
        10'd 147:out = 12'd 1552;
        10'd 148:out = 12'd 1557;
        10'd 149:out = 12'd 1562;
        10'd 150:out = 12'd 1568;
        10'd 151:out = 12'd 1573;
        10'd 152:out = 12'd 1578;
        10'd 153:out = 12'd 1583;
        10'd 154:out = 12'd 1588;
        10'd 155:out = 12'd 1594;
        10'd 156:out = 12'd 1599;
        10'd 157:out = 12'd 1604;
        10'd 158:out = 12'd 1609;
        10'd 159:out = 12'd 1614;
        10'd 160:out = 12'd 1619;
        10'd 161:out = 12'd 1624;
        10'd 162:out = 12'd 1629;
        10'd 163:out = 12'd 1634;
        10'd 164:out = 12'd 1639;
        10'd 165:out = 12'd 1644;
        10'd 166:out = 12'd 1649;
        10'd 167:out = 12'd 1654;
        10'd 168:out = 12'd 1659;
        10'd 169:out = 12'd 1664;
        10'd 170:out = 12'd 1669;
        10'd 171:out = 12'd 1674;
        10'd 172:out = 12'd 1679;
        10'd 173:out = 12'd 1684;
        10'd 174:out = 12'd 1688;
        10'd 175:out = 12'd 1693;
        10'd 176:out = 12'd 1698;
        10'd 177:out = 12'd 1703;
        10'd 178:out = 12'd 1708;
        10'd 179:out = 12'd 1713;
        10'd 180:out = 12'd 1717;
        10'd 181:out = 12'd 1722;
        10'd 182:out = 12'd 1727;
        10'd 183:out = 12'd 1732;
        10'd 184:out = 12'd 1736;
        10'd 185:out = 12'd 1741;
        10'd 186:out = 12'd 1746;
        10'd 187:out = 12'd 1750;
        10'd 188:out = 12'd 1755;
        10'd 189:out = 12'd 1760;
        10'd 190:out = 12'd 1764;
        10'd 191:out = 12'd 1769;
        10'd 192:out = 12'd 1774;
        10'd 193:out = 12'd 1778;
        10'd 194:out = 12'd 1783;
        10'd 195:out = 12'd 1787;
        10'd 196:out = 12'd 1792;
        10'd 197:out = 12'd 1797;
        10'd 198:out = 12'd 1801;
        10'd 199:out = 12'd 1806;
        10'd 200:out = 12'd 1810;
        10'd 201:out = 12'd 1815;
        10'd 202:out = 12'd 1819;
        10'd 203:out = 12'd 1824;
        10'd 204:out = 12'd 1828;
        10'd 205:out = 12'd 1833;
        10'd 206:out = 12'd 1837;
        10'd 207:out = 12'd 1842;
        10'd 208:out = 12'd 1846;
        10'd 209:out = 12'd 1850;
        10'd 210:out = 12'd 1855;
        10'd 211:out = 12'd 1859;
        10'd 212:out = 12'd 1864;
        10'd 213:out = 12'd 1868;
        10'd 214:out = 12'd 1872;
        10'd 215:out = 12'd 1877;
        10'd 216:out = 12'd 1881;
        10'd 217:out = 12'd 1886;
        10'd 218:out = 12'd 1890;
        10'd 219:out = 12'd 1894;
        10'd 220:out = 12'd 1899;
        10'd 221:out = 12'd 1903;
        10'd 222:out = 12'd 1907;
        10'd 223:out = 12'd 1911;
        10'd 224:out = 12'd 1916;
        10'd 225:out = 12'd 1920;
        10'd 226:out = 12'd 1924;
        10'd 227:out = 12'd 1929;
        10'd 228:out = 12'd 1933;
        10'd 229:out = 12'd 1937;
        10'd 230:out = 12'd 1941;
        10'd 231:out = 12'd 1945;
        10'd 232:out = 12'd 1950;
        10'd 233:out = 12'd 1954;
        10'd 234:out = 12'd 1958;
        10'd 235:out = 12'd 1962;
        10'd 236:out = 12'd 1966;
        10'd 237:out = 12'd 1971;
        10'd 238:out = 12'd 1975;
        10'd 239:out = 12'd 1979;
        10'd 240:out = 12'd 1983;
        10'd 241:out = 12'd 1987;
        10'd 242:out = 12'd 1991;
        10'd 243:out = 12'd 1995;
        10'd 244:out = 12'd 1999;
        10'd 245:out = 12'd 2004;
        10'd 246:out = 12'd 2008;
        10'd 247:out = 12'd 2012;
        10'd 248:out = 12'd 2016;
        10'd 249:out = 12'd 2020;
        10'd 250:out = 12'd 2024;
        10'd 251:out = 12'd 2028;
        10'd 252:out = 12'd 2032;
        10'd 253:out = 12'd 2036;
        10'd 254:out = 12'd 2040;
        10'd 255:out = 12'd 2044;
        10'd 256:out = 12'd 2048;
        10'd 257:out = 12'd 2052;
        10'd 258:out = 12'd 2056;
        10'd 259:out = 12'd 2060;
        10'd 260:out = 12'd 2064;
        10'd 261:out = 12'd 2068;
        10'd 262:out = 12'd 2072;
        10'd 263:out = 12'd 2076;
        10'd 264:out = 12'd 2080;
        10'd 265:out = 12'd 2084;
        10'd 266:out = 12'd 2088;
        10'd 267:out = 12'd 2092;
        10'd 268:out = 12'd 2095;
        10'd 269:out = 12'd 2099;
        10'd 270:out = 12'd 2103;
        10'd 271:out = 12'd 2107;
        10'd 272:out = 12'd 2111;
        10'd 273:out = 12'd 2115;
        10'd 274:out = 12'd 2119;
        10'd 275:out = 12'd 2123;
        10'd 276:out = 12'd 2126;
        10'd 277:out = 12'd 2130;
        10'd 278:out = 12'd 2134;
        10'd 279:out = 12'd 2138;
        10'd 280:out = 12'd 2142;
        10'd 281:out = 12'd 2146;
        10'd 282:out = 12'd 2149;
        10'd 283:out = 12'd 2153;
        10'd 284:out = 12'd 2157;
        10'd 285:out = 12'd 2161;
        10'd 286:out = 12'd 2165;
        10'd 287:out = 12'd 2168;
        10'd 288:out = 12'd 2172;
        10'd 289:out = 12'd 2176;
        10'd 290:out = 12'd 2180;
        10'd 291:out = 12'd 2184;
        10'd 292:out = 12'd 2187;
        10'd 293:out = 12'd 2191;
        10'd 294:out = 12'd 2195;
        10'd 295:out = 12'd 2198;
        10'd 296:out = 12'd 2202;
        10'd 297:out = 12'd 2206;
        10'd 298:out = 12'd 2210;
        10'd 299:out = 12'd 2213;
        10'd 300:out = 12'd 2217;
        10'd 301:out = 12'd 2221;
        10'd 302:out = 12'd 2224;
        10'd 303:out = 12'd 2228;
        10'd 304:out = 12'd 2232;
        10'd 305:out = 12'd 2235;
        10'd 306:out = 12'd 2239;
        10'd 307:out = 12'd 2243;
        10'd 308:out = 12'd 2246;
        10'd 309:out = 12'd 2250;
        10'd 310:out = 12'd 2254;
        10'd 311:out = 12'd 2257;
        10'd 312:out = 12'd 2261;
        10'd 313:out = 12'd 2265;
        10'd 314:out = 12'd 2268;
        10'd 315:out = 12'd 2272;
        10'd 316:out = 12'd 2275;
        10'd 317:out = 12'd 2279;
        10'd 318:out = 12'd 2283;
        10'd 319:out = 12'd 2286;
        10'd 320:out = 12'd 2290;
        10'd 321:out = 12'd 2293;
        10'd 322:out = 12'd 2297;
        10'd 323:out = 12'd 2300;
        10'd 324:out = 12'd 2304;
        10'd 325:out = 12'd 2308;
        10'd 326:out = 12'd 2311;
        10'd 327:out = 12'd 2315;
        10'd 328:out = 12'd 2318;
        10'd 329:out = 12'd 2322;
        10'd 330:out = 12'd 2325;
        10'd 331:out = 12'd 2329;
        10'd 332:out = 12'd 2332;
        10'd 333:out = 12'd 2336;
        10'd 334:out = 12'd 2339;
        10'd 335:out = 12'd 2343;
        10'd 336:out = 12'd 2346;
        10'd 337:out = 12'd 2350;
        10'd 338:out = 12'd 2353;
        10'd 339:out = 12'd 2357;
        10'd 340:out = 12'd 2360;
        10'd 341:out = 12'd 2364;
        10'd 342:out = 12'd 2367;
        10'd 343:out = 12'd 2371;
        10'd 344:out = 12'd 2374;
        10'd 345:out = 12'd 2377;
        10'd 346:out = 12'd 2381;
        10'd 347:out = 12'd 2384;
        10'd 348:out = 12'd 2388;
        10'd 349:out = 12'd 2391;
        10'd 350:out = 12'd 2395;
        10'd 351:out = 12'd 2398;
        10'd 352:out = 12'd 2401;
        10'd 353:out = 12'd 2405;
        10'd 354:out = 12'd 2408;
        10'd 355:out = 12'd 2412;
        10'd 356:out = 12'd 2415;
        10'd 357:out = 12'd 2418;
        10'd 358:out = 12'd 2422;
        10'd 359:out = 12'd 2425;
        10'd 360:out = 12'd 2429;
        10'd 361:out = 12'd 2432;
        10'd 362:out = 12'd 2435;
        10'd 363:out = 12'd 2439;
        10'd 364:out = 12'd 2442;
        10'd 365:out = 12'd 2445;
        10'd 366:out = 12'd 2449;
        10'd 367:out = 12'd 2452;
        10'd 368:out = 12'd 2455;
        10'd 369:out = 12'd 2459;
        10'd 370:out = 12'd 2462;
        10'd 371:out = 12'd 2465;
        10'd 372:out = 12'd 2469;
        10'd 373:out = 12'd 2472;
        10'd 374:out = 12'd 2475;
        10'd 375:out = 12'd 2479;
        10'd 376:out = 12'd 2482;
        10'd 377:out = 12'd 2485;
        10'd 378:out = 12'd 2489;
        10'd 379:out = 12'd 2492;
        10'd 380:out = 12'd 2495;
        10'd 381:out = 12'd 2498;
        10'd 382:out = 12'd 2502;
        10'd 383:out = 12'd 2505;
        10'd 384:out = 12'd 2508;
        10'd 385:out = 12'd 2512;
        10'd 386:out = 12'd 2515;
        10'd 387:out = 12'd 2518;
        10'd 388:out = 12'd 2521;
        10'd 389:out = 12'd 2525;
        10'd 390:out = 12'd 2528;
        10'd 391:out = 12'd 2531;
        10'd 392:out = 12'd 2534;
        10'd 393:out = 12'd 2538;
        10'd 394:out = 12'd 2541;
        10'd 395:out = 12'd 2544;
        10'd 396:out = 12'd 2547;
        10'd 397:out = 12'd 2550;
        10'd 398:out = 12'd 2554;
        10'd 399:out = 12'd 2557;
        10'd 400:out = 12'd 2560;
        10'd 401:out = 12'd 2563;
        10'd 402:out = 12'd 2566;
        10'd 403:out = 12'd 2570;
        10'd 404:out = 12'd 2573;
        10'd 405:out = 12'd 2576;
        10'd 406:out = 12'd 2579;
        10'd 407:out = 12'd 2582;
        10'd 408:out = 12'd 2585;
        10'd 409:out = 12'd 2589;
        10'd 410:out = 12'd 2592;
        10'd 411:out = 12'd 2595;
        10'd 412:out = 12'd 2598;
        10'd 413:out = 12'd 2601;
        10'd 414:out = 12'd 2604;
        10'd 415:out = 12'd 2608;
        10'd 416:out = 12'd 2611;
        10'd 417:out = 12'd 2614;
        10'd 418:out = 12'd 2617;
        10'd 419:out = 12'd 2620;
        10'd 420:out = 12'd 2623;
        10'd 421:out = 12'd 2626;
        10'd 422:out = 12'd 2629;
        10'd 423:out = 12'd 2633;
        10'd 424:out = 12'd 2636;
        10'd 425:out = 12'd 2639;
        10'd 426:out = 12'd 2642;
        10'd 427:out = 12'd 2645;
        10'd 428:out = 12'd 2648;
        10'd 429:out = 12'd 2651;
        10'd 430:out = 12'd 2654;
        10'd 431:out = 12'd 2657;
        10'd 432:out = 12'd 2660;
        10'd 433:out = 12'd 2664;
        10'd 434:out = 12'd 2667;
        10'd 435:out = 12'd 2670;
        10'd 436:out = 12'd 2673;
        10'd 437:out = 12'd 2676;
        10'd 438:out = 12'd 2679;
        10'd 439:out = 12'd 2682;
        10'd 440:out = 12'd 2685;
        10'd 441:out = 12'd 2688;
        10'd 442:out = 12'd 2691;
        10'd 443:out = 12'd 2694;
        10'd 444:out = 12'd 2697;
        10'd 445:out = 12'd 2700;
        10'd 446:out = 12'd 2703;
        10'd 447:out = 12'd 2706;
        10'd 448:out = 12'd 2709;
        10'd 449:out = 12'd 2712;
        10'd 450:out = 12'd 2715;
        10'd 451:out = 12'd 2718;
        10'd 452:out = 12'd 2721;
        10'd 453:out = 12'd 2724;
        10'd 454:out = 12'd 2727;
        10'd 455:out = 12'd 2730;
        10'd 456:out = 12'd 2733;
        10'd 457:out = 12'd 2736;
        10'd 458:out = 12'd 2739;
        10'd 459:out = 12'd 2742;
        10'd 460:out = 12'd 2745;
        10'd 461:out = 12'd 2748;
        10'd 462:out = 12'd 2751;
        10'd 463:out = 12'd 2754;
        10'd 464:out = 12'd 2757;
        10'd 465:out = 12'd 2760;
        10'd 466:out = 12'd 2763;
        10'd 467:out = 12'd 2766;
        10'd 468:out = 12'd 2769;
        10'd 469:out = 12'd 2772;
        10'd 470:out = 12'd 2775;
        10'd 471:out = 12'd 2778;
        10'd 472:out = 12'd 2781;
        10'd 473:out = 12'd 2784;
        10'd 474:out = 12'd 2787;
        10'd 475:out = 12'd 2790;
        10'd 476:out = 12'd 2793;
        10'd 477:out = 12'd 2796;
        10'd 478:out = 12'd 2798;
        10'd 479:out = 12'd 2801;
        10'd 480:out = 12'd 2804;
        10'd 481:out = 12'd 2807;
        10'd 482:out = 12'd 2810;
        10'd 483:out = 12'd 2813;
        10'd 484:out = 12'd 2816;
        10'd 485:out = 12'd 2819;
        10'd 486:out = 12'd 2822;
        10'd 487:out = 12'd 2825;
        10'd 488:out = 12'd 2828;
        10'd 489:out = 12'd 2831;
        10'd 490:out = 12'd 2833;
        10'd 491:out = 12'd 2836;
        10'd 492:out = 12'd 2839;
        10'd 493:out = 12'd 2842;
        10'd 494:out = 12'd 2845;
        10'd 495:out = 12'd 2848;
        10'd 496:out = 12'd 2851;
        10'd 497:out = 12'd 2854;
        10'd 498:out = 12'd 2856;
        10'd 499:out = 12'd 2859;
        10'd 500:out = 12'd 2862;
        10'd 501:out = 12'd 2865;
        10'd 502:out = 12'd 2868;
        10'd 503:out = 12'd 2871;
        10'd 504:out = 12'd 2874;
        10'd 505:out = 12'd 2876;
        10'd 506:out = 12'd 2879;
        10'd 507:out = 12'd 2882;
        10'd 508:out = 12'd 2885;
        10'd 509:out = 12'd 2888;
        10'd 510:out = 12'd 2891;
        10'd 511:out = 12'd 2893;
        10'd 512:out = 12'd 2896;
        10'd 513:out = 12'd 2899;
        10'd 514:out = 12'd 2902;
        10'd 515:out = 12'd 2905;
        10'd 516:out = 12'd 2908;
        10'd 517:out = 12'd 2910;
        10'd 518:out = 12'd 2913;
        10'd 519:out = 12'd 2916;
        10'd 520:out = 12'd 2919;
        10'd 521:out = 12'd 2922;
        10'd 522:out = 12'd 2924;
        10'd 523:out = 12'd 2927;
        10'd 524:out = 12'd 2930;
        10'd 525:out = 12'd 2933;
        10'd 526:out = 12'd 2936;
        10'd 527:out = 12'd 2938;
        10'd 528:out = 12'd 2941;
        10'd 529:out = 12'd 2944;
        10'd 530:out = 12'd 2947;
        10'd 531:out = 12'd 2950;
        10'd 532:out = 12'd 2952;
        10'd 533:out = 12'd 2955;
        10'd 534:out = 12'd 2958;
        10'd 535:out = 12'd 2961;
        10'd 536:out = 12'd 2963;
        10'd 537:out = 12'd 2966;
        10'd 538:out = 12'd 2969;
        10'd 539:out = 12'd 2972;
        10'd 540:out = 12'd 2974;
        10'd 541:out = 12'd 2977;
        10'd 542:out = 12'd 2980;
        10'd 543:out = 12'd 2983;
        10'd 544:out = 12'd 2985;
        10'd 545:out = 12'd 2988;
        10'd 546:out = 12'd 2991;
        10'd 547:out = 12'd 2994;
        10'd 548:out = 12'd 2996;
        10'd 549:out = 12'd 2999;
        10'd 550:out = 12'd 3002;
        10'd 551:out = 12'd 3005;
        10'd 552:out = 12'd 3007;
        10'd 553:out = 12'd 3010;
        10'd 554:out = 12'd 3013;
        10'd 555:out = 12'd 3015;
        10'd 556:out = 12'd 3018;
        10'd 557:out = 12'd 3021;
        10'd 558:out = 12'd 3024;
        10'd 559:out = 12'd 3026;
        10'd 560:out = 12'd 3029;
        10'd 561:out = 12'd 3032;
        10'd 562:out = 12'd 3034;
        10'd 563:out = 12'd 3037;
        10'd 564:out = 12'd 3040;
        10'd 565:out = 12'd 3043;
        10'd 566:out = 12'd 3045;
        10'd 567:out = 12'd 3048;
        10'd 568:out = 12'd 3051;
        10'd 569:out = 12'd 3053;
        10'd 570:out = 12'd 3056;
        10'd 571:out = 12'd 3059;
        10'd 572:out = 12'd 3061;
        10'd 573:out = 12'd 3064;
        10'd 574:out = 12'd 3067;
        10'd 575:out = 12'd 3069;
        10'd 576:out = 12'd 3072;
        10'd 577:out = 12'd 3075;
        10'd 578:out = 12'd 3077;
        10'd 579:out = 12'd 3080;
        10'd 580:out = 12'd 3083;
        10'd 581:out = 12'd 3085;
        10'd 582:out = 12'd 3088;
        10'd 583:out = 12'd 3091;
        10'd 584:out = 12'd 3093;
        10'd 585:out = 12'd 3096;
        10'd 586:out = 12'd 3099;
        10'd 587:out = 12'd 3101;
        10'd 588:out = 12'd 3104;
        10'd 589:out = 12'd 3106;
        10'd 590:out = 12'd 3109;
        10'd 591:out = 12'd 3112;
        10'd 592:out = 12'd 3114;
        10'd 593:out = 12'd 3117;
        10'd 594:out = 12'd 3120;
        10'd 595:out = 12'd 3122;
        10'd 596:out = 12'd 3125;
        10'd 597:out = 12'd 3127;
        10'd 598:out = 12'd 3130;
        10'd 599:out = 12'd 3133;
        10'd 600:out = 12'd 3135;
        10'd 601:out = 12'd 3138;
        10'd 602:out = 12'd 3141;
        10'd 603:out = 12'd 3143;
        10'd 604:out = 12'd 3146;
        10'd 605:out = 12'd 3148;
        10'd 606:out = 12'd 3151;
        10'd 607:out = 12'd 3154;
        10'd 608:out = 12'd 3156;
        10'd 609:out = 12'd 3159;
        10'd 610:out = 12'd 3161;
        10'd 611:out = 12'd 3164;
        10'd 612:out = 12'd 3167;
        10'd 613:out = 12'd 3169;
        10'd 614:out = 12'd 3172;
        10'd 615:out = 12'd 3174;
        10'd 616:out = 12'd 3177;
        10'd 617:out = 12'd 3179;
        10'd 618:out = 12'd 3182;
        10'd 619:out = 12'd 3185;
        10'd 620:out = 12'd 3187;
        10'd 621:out = 12'd 3190;
        10'd 622:out = 12'd 3192;
        10'd 623:out = 12'd 3195;
        10'd 624:out = 12'd 3197;
        10'd 625:out = 12'd 3200;
        10'd 626:out = 12'd 3203;
        10'd 627:out = 12'd 3205;
        10'd 628:out = 12'd 3208;
        10'd 629:out = 12'd 3210;
        10'd 630:out = 12'd 3213;
        10'd 631:out = 12'd 3215;
        10'd 632:out = 12'd 3218;
        10'd 633:out = 12'd 3220;
        10'd 634:out = 12'd 3223;
        10'd 635:out = 12'd 3225;
        10'd 636:out = 12'd 3228;
        10'd 637:out = 12'd 3231;
        10'd 638:out = 12'd 3233;
        10'd 639:out = 12'd 3236;
        10'd 640:out = 12'd 3238;
        10'd 641:out = 12'd 3241;
        10'd 642:out = 12'd 3243;
        10'd 643:out = 12'd 3246;
        10'd 644:out = 12'd 3248;
        10'd 645:out = 12'd 3251;
        10'd 646:out = 12'd 3253;
        10'd 647:out = 12'd 3256;
        10'd 648:out = 12'd 3258;
        10'd 649:out = 12'd 3261;
        10'd 650:out = 12'd 3263;
        10'd 651:out = 12'd 3266;
        10'd 652:out = 12'd 3268;
        10'd 653:out = 12'd 3271;
        10'd 654:out = 12'd 3273;
        10'd 655:out = 12'd 3276;
        10'd 656:out = 12'd 3278;
        10'd 657:out = 12'd 3281;
        10'd 658:out = 12'd 3283;
        10'd 659:out = 12'd 3286;
        10'd 660:out = 12'd 3288;
        10'd 661:out = 12'd 3291;
        10'd 662:out = 12'd 3293;
        10'd 663:out = 12'd 3296;
        10'd 664:out = 12'd 3298;
        10'd 665:out = 12'd 3301;
        10'd 666:out = 12'd 3303;
        10'd 667:out = 12'd 3306;
        10'd 668:out = 12'd 3308;
        10'd 669:out = 12'd 3311;
        10'd 670:out = 12'd 3313;
        10'd 671:out = 12'd 3316;
        10'd 672:out = 12'd 3318;
        10'd 673:out = 12'd 3321;
        10'd 674:out = 12'd 3323;
        10'd 675:out = 12'd 3326;
        10'd 676:out = 12'd 3328;
        10'd 677:out = 12'd 3330;
        10'd 678:out = 12'd 3333;
        10'd 679:out = 12'd 3335;
        10'd 680:out = 12'd 3338;
        10'd 681:out = 12'd 3340;
        10'd 682:out = 12'd 3343;
        10'd 683:out = 12'd 3345;
        10'd 684:out = 12'd 3348;
        10'd 685:out = 12'd 3350;
        10'd 686:out = 12'd 3353;
        10'd 687:out = 12'd 3355;
        10'd 688:out = 12'd 3357;
        10'd 689:out = 12'd 3360;
        10'd 690:out = 12'd 3362;
        10'd 691:out = 12'd 3365;
        10'd 692:out = 12'd 3367;
        10'd 693:out = 12'd 3370;
        10'd 694:out = 12'd 3372;
        10'd 695:out = 12'd 3374;
        10'd 696:out = 12'd 3377;
        10'd 697:out = 12'd 3379;
        10'd 698:out = 12'd 3382;
        10'd 699:out = 12'd 3384;
        10'd 700:out = 12'd 3387;
        10'd 701:out = 12'd 3389;
        10'd 702:out = 12'd 3391;
        10'd 703:out = 12'd 3394;
        10'd 704:out = 12'd 3396;
        10'd 705:out = 12'd 3399;
        10'd 706:out = 12'd 3401;
        10'd 707:out = 12'd 3403;
        10'd 708:out = 12'd 3406;
        10'd 709:out = 12'd 3408;
        10'd 710:out = 12'd 3411;
        10'd 711:out = 12'd 3413;
        10'd 712:out = 12'd 3415;
        10'd 713:out = 12'd 3418;
        10'd 714:out = 12'd 3420;
        10'd 715:out = 12'd 3423;
        10'd 716:out = 12'd 3425;
        10'd 717:out = 12'd 3427;
        10'd 718:out = 12'd 3430;
        10'd 719:out = 12'd 3432;
        10'd 720:out = 12'd 3435;
        10'd 721:out = 12'd 3437;
        10'd 722:out = 12'd 3439;
        10'd 723:out = 12'd 3442;
        10'd 724:out = 12'd 3444;
        10'd 725:out = 12'd 3447;
        10'd 726:out = 12'd 3449;
        10'd 727:out = 12'd 3451;
        10'd 728:out = 12'd 3454;
        10'd 729:out = 12'd 3456;
        10'd 730:out = 12'd 3458;
        10'd 731:out = 12'd 3461;
        10'd 732:out = 12'd 3463;
        10'd 733:out = 12'd 3465;
        10'd 734:out = 12'd 3468;
        10'd 735:out = 12'd 3470;
        10'd 736:out = 12'd 3473;
        10'd 737:out = 12'd 3475;
        10'd 738:out = 12'd 3477;
        10'd 739:out = 12'd 3480;
        10'd 740:out = 12'd 3482;
        10'd 741:out = 12'd 3484;
        10'd 742:out = 12'd 3487;
        10'd 743:out = 12'd 3489;
        10'd 744:out = 12'd 3491;
        10'd 745:out = 12'd 3494;
        10'd 746:out = 12'd 3496;
        10'd 747:out = 12'd 3498;
        10'd 748:out = 12'd 3501;
        10'd 749:out = 12'd 3503;
        10'd 750:out = 12'd 3505;
        10'd 751:out = 12'd 3508;
        10'd 752:out = 12'd 3510;
        10'd 753:out = 12'd 3512;
        10'd 754:out = 12'd 3515;
        10'd 755:out = 12'd 3517;
        10'd 756:out = 12'd 3519;
        10'd 757:out = 12'd 3522;
        10'd 758:out = 12'd 3524;
        10'd 759:out = 12'd 3526;
        10'd 760:out = 12'd 3529;
        10'd 761:out = 12'd 3531;
        10'd 762:out = 12'd 3533;
        10'd 763:out = 12'd 3536;
        10'd 764:out = 12'd 3538;
        10'd 765:out = 12'd 3540;
        10'd 766:out = 12'd 3543;
        10'd 767:out = 12'd 3545;
        10'd 768:out = 12'd 3547;
        10'd 769:out = 12'd 3550;
        10'd 770:out = 12'd 3552;
        10'd 771:out = 12'd 3554;
        10'd 772:out = 12'd 3556;
        10'd 773:out = 12'd 3559;
        10'd 774:out = 12'd 3561;
        10'd 775:out = 12'd 3563;
        10'd 776:out = 12'd 3566;
        10'd 777:out = 12'd 3568;
        10'd 778:out = 12'd 3570;
        10'd 779:out = 12'd 3573;
        10'd 780:out = 12'd 3575;
        10'd 781:out = 12'd 3577;
        10'd 782:out = 12'd 3579;
        10'd 783:out = 12'd 3582;
        10'd 784:out = 12'd 3584;
        10'd 785:out = 12'd 3586;
        10'd 786:out = 12'd 3589;
        10'd 787:out = 12'd 3591;
        10'd 788:out = 12'd 3593;
        10'd 789:out = 12'd 3595;
        10'd 790:out = 12'd 3598;
        10'd 791:out = 12'd 3600;
        10'd 792:out = 12'd 3602;
        10'd 793:out = 12'd 3605;
        10'd 794:out = 12'd 3607;
        10'd 795:out = 12'd 3609;
        10'd 796:out = 12'd 3611;
        10'd 797:out = 12'd 3614;
        10'd 798:out = 12'd 3616;
        10'd 799:out = 12'd 3618;
        10'd 800:out = 12'd 3620;
        10'd 801:out = 12'd 3623;
        10'd 802:out = 12'd 3625;
        10'd 803:out = 12'd 3627;
        10'd 804:out = 12'd 3629;
        10'd 805:out = 12'd 3632;
        10'd 806:out = 12'd 3634;
        10'd 807:out = 12'd 3636;
        10'd 808:out = 12'd 3638;
        10'd 809:out = 12'd 3641;
        10'd 810:out = 12'd 3643;
        10'd 811:out = 12'd 3645;
        10'd 812:out = 12'd 3647;
        10'd 813:out = 12'd 3650;
        10'd 814:out = 12'd 3652;
        10'd 815:out = 12'd 3654;
        10'd 816:out = 12'd 3656;
        10'd 817:out = 12'd 3659;
        10'd 818:out = 12'd 3661;
        10'd 819:out = 12'd 3663;
        10'd 820:out = 12'd 3665;
        10'd 821:out = 12'd 3668;
        10'd 822:out = 12'd 3670;
        10'd 823:out = 12'd 3672;
        10'd 824:out = 12'd 3674;
        10'd 825:out = 12'd 3677;
        10'd 826:out = 12'd 3679;
        10'd 827:out = 12'd 3681;
        10'd 828:out = 12'd 3683;
        10'd 829:out = 12'd 3685;
        10'd 830:out = 12'd 3688;
        10'd 831:out = 12'd 3690;
        10'd 832:out = 12'd 3692;
        10'd 833:out = 12'd 3694;
        10'd 834:out = 12'd 3697;
        10'd 835:out = 12'd 3699;
        10'd 836:out = 12'd 3701;
        10'd 837:out = 12'd 3703;
        10'd 838:out = 12'd 3705;
        10'd 839:out = 12'd 3708;
        10'd 840:out = 12'd 3710;
        10'd 841:out = 12'd 3712;
        10'd 842:out = 12'd 3714;
        10'd 843:out = 12'd 3716;
        10'd 844:out = 12'd 3719;
        10'd 845:out = 12'd 3721;
        10'd 846:out = 12'd 3723;
        10'd 847:out = 12'd 3725;
        10'd 848:out = 12'd 3727;
        10'd 849:out = 12'd 3730;
        10'd 850:out = 12'd 3732;
        10'd 851:out = 12'd 3734;
        10'd 852:out = 12'd 3736;
        10'd 853:out = 12'd 3738;
        10'd 854:out = 12'd 3741;
        10'd 855:out = 12'd 3743;
        10'd 856:out = 12'd 3745;
        10'd 857:out = 12'd 3747;
        10'd 858:out = 12'd 3749;
        10'd 859:out = 12'd 3752;
        10'd 860:out = 12'd 3754;
        10'd 861:out = 12'd 3756;
        10'd 862:out = 12'd 3758;
        10'd 863:out = 12'd 3760;
        10'd 864:out = 12'd 3762;
        10'd 865:out = 12'd 3765;
        10'd 866:out = 12'd 3767;
        10'd 867:out = 12'd 3769;
        10'd 868:out = 12'd 3771;
        10'd 869:out = 12'd 3773;
        10'd 870:out = 12'd 3775;
        10'd 871:out = 12'd 3778;
        10'd 872:out = 12'd 3780;
        10'd 873:out = 12'd 3782;
        10'd 874:out = 12'd 3784;
        10'd 875:out = 12'd 3786;
        10'd 876:out = 12'd 3788;
        10'd 877:out = 12'd 3791;
        10'd 878:out = 12'd 3793;
        10'd 879:out = 12'd 3795;
        10'd 880:out = 12'd 3797;
        10'd 881:out = 12'd 3799;
        10'd 882:out = 12'd 3801;
        10'd 883:out = 12'd 3804;
        10'd 884:out = 12'd 3806;
        10'd 885:out = 12'd 3808;
        10'd 886:out = 12'd 3810;
        10'd 887:out = 12'd 3812;
        10'd 888:out = 12'd 3814;
        10'd 889:out = 12'd 3816;
        10'd 890:out = 12'd 3819;
        10'd 891:out = 12'd 3821;
        10'd 892:out = 12'd 3823;
        10'd 893:out = 12'd 3825;
        10'd 894:out = 12'd 3827;
        10'd 895:out = 12'd 3829;
        10'd 896:out = 12'd 3831;
        10'd 897:out = 12'd 3834;
        10'd 898:out = 12'd 3836;
        10'd 899:out = 12'd 3838;
        10'd 900:out = 12'd 3840;
        10'd 901:out = 12'd 3842;
        10'd 902:out = 12'd 3844;
        10'd 903:out = 12'd 3846;
        10'd 904:out = 12'd 3849;
        10'd 905:out = 12'd 3851;
        10'd 906:out = 12'd 3853;
        10'd 907:out = 12'd 3855;
        10'd 908:out = 12'd 3857;
        10'd 909:out = 12'd 3859;
        10'd 910:out = 12'd 3861;
        10'd 911:out = 12'd 3863;
        10'd 912:out = 12'd 3866;
        10'd 913:out = 12'd 3868;
        10'd 914:out = 12'd 3870;
        10'd 915:out = 12'd 3872;
        10'd 916:out = 12'd 3874;
        10'd 917:out = 12'd 3876;
        10'd 918:out = 12'd 3878;
        10'd 919:out = 12'd 3880;
        10'd 920:out = 12'd 3882;
        10'd 921:out = 12'd 3885;
        10'd 922:out = 12'd 3887;
        10'd 923:out = 12'd 3889;
        10'd 924:out = 12'd 3891;
        10'd 925:out = 12'd 3893;
        10'd 926:out = 12'd 3895;
        10'd 927:out = 12'd 3897;
        10'd 928:out = 12'd 3899;
        10'd 929:out = 12'd 3901;
        10'd 930:out = 12'd 3903;
        10'd 931:out = 12'd 3906;
        10'd 932:out = 12'd 3908;
        10'd 933:out = 12'd 3910;
        10'd 934:out = 12'd 3912;
        10'd 935:out = 12'd 3914;
        10'd 936:out = 12'd 3916;
        10'd 937:out = 12'd 3918;
        10'd 938:out = 12'd 3920;
        10'd 939:out = 12'd 3922;
        10'd 940:out = 12'd 3924;
        10'd 941:out = 12'd 3926;
        10'd 942:out = 12'd 3929;
        10'd 943:out = 12'd 3931;
        10'd 944:out = 12'd 3933;
        10'd 945:out = 12'd 3935;
        10'd 946:out = 12'd 3937;
        10'd 947:out = 12'd 3939;
        10'd 948:out = 12'd 3941;
        10'd 949:out = 12'd 3943;
        10'd 950:out = 12'd 3945;
        10'd 951:out = 12'd 3947;
        10'd 952:out = 12'd 3949;
        10'd 953:out = 12'd 3951;
        10'd 954:out = 12'd 3954;
        10'd 955:out = 12'd 3956;
        10'd 956:out = 12'd 3958;
        10'd 957:out = 12'd 3960;
        10'd 958:out = 12'd 3962;
        10'd 959:out = 12'd 3964;
        10'd 960:out = 12'd 3966;
        10'd 961:out = 12'd 3968;
        10'd 962:out = 12'd 3970;
        10'd 963:out = 12'd 3972;
        10'd 964:out = 12'd 3974;
        10'd 965:out = 12'd 3976;
        10'd 966:out = 12'd 3978;
        10'd 967:out = 12'd 3980;
        10'd 968:out = 12'd 3982;
        10'd 969:out = 12'd 3984;
        10'd 970:out = 12'd 3987;
        10'd 971:out = 12'd 3989;
        10'd 972:out = 12'd 3991;
        10'd 973:out = 12'd 3993;
        10'd 974:out = 12'd 3995;
        10'd 975:out = 12'd 3997;
        10'd 976:out = 12'd 3999;
        10'd 977:out = 12'd 4001;
        10'd 978:out = 12'd 4003;
        10'd 979:out = 12'd 4005;
        10'd 980:out = 12'd 4007;
        10'd 981:out = 12'd 4009;
        10'd 982:out = 12'd 4011;
        10'd 983:out = 12'd 4013;
        10'd 984:out = 12'd 4015;
        10'd 985:out = 12'd 4017;
        10'd 986:out = 12'd 4019;
        10'd 987:out = 12'd 4021;
        10'd 988:out = 12'd 4023;
        10'd 989:out = 12'd 4025;
        10'd 990:out = 12'd 4027;
        10'd 991:out = 12'd 4029;
        10'd 992:out = 12'd 4031;
        10'd 993:out = 12'd 4034;
        10'd 994:out = 12'd 4036;
        10'd 995:out = 12'd 4038;
        10'd 996:out = 12'd 4040;
        10'd 997:out = 12'd 4042;
        10'd 998:out = 12'd 4044;
        10'd 999:out = 12'd 4046;
        10'd 1000:out = 12'd 4048;
        10'd 1001:out = 12'd 4050;
        10'd 1002:out = 12'd 4052;
        10'd 1003:out = 12'd 4054;
        10'd 1004:out = 12'd 4056;
        10'd 1005:out = 12'd 4058;
        10'd 1006:out = 12'd 4060;
        10'd 1007:out = 12'd 4062;
        10'd 1008:out = 12'd 4064;
        10'd 1009:out = 12'd 4066;
        10'd 1010:out = 12'd 4068;
        10'd 1011:out = 12'd 4070;
        10'd 1012:out = 12'd 4072;
        10'd 1013:out = 12'd 4074;
        10'd 1014:out = 12'd 4076;
        10'd 1015:out = 12'd 4078;
        10'd 1016:out = 12'd 4080;
        10'd 1017:out = 12'd 4082;
        10'd 1018:out = 12'd 4084;
        10'd 1019:out = 12'd 4086;
        10'd 1020:out = 12'd 4088;
        10'd 1021:out = 12'd 4090;
        10'd 1022:out = 12'd 4092;
        10'd 1023:out = 12'd 4094;
            default:    out = 12'd0;
        endcase
    end    
    
endmodule
