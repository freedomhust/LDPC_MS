/*
 * Author: neidong_fu
 * Time  : 2020/03/04
 * function: caculate cos(x)
*/

module cos_quad_LUT(
    // out = ceil((2^14-1)*cos(2*pi*in/2^12))
    input [10:0] in,
    output reg [13:0] out
    );
    
    always@(*) begin
        case(in)
            11'd 1:out = 14'd 16383;
        11'd 2:out = 14'd 16383;
        11'd 3:out = 14'd 16383;
        11'd 4:out = 14'd 16383;
        11'd 5:out = 14'd 16383;
        11'd 6:out = 14'd 16383;
        11'd 7:out = 14'd 16383;
        11'd 8:out = 14'd 16382;
        11'd 9:out = 14'd 16382;
        11'd 10:out = 14'd 16382;
        11'd 11:out = 14'd 16381;
        11'd 12:out = 14'd 16381;
        11'd 13:out = 14'd 16380;
        11'd 14:out = 14'd 16380;
        11'd 15:out = 14'd 16379;
        11'd 16:out = 14'd 16379;
        11'd 17:out = 14'd 16378;
        11'd 18:out = 14'd 16377;
        11'd 19:out = 14'd 16377;
        11'd 20:out = 14'd 16376;
        11'd 21:out = 14'd 16375;
        11'd 22:out = 14'd 16374;
        11'd 23:out = 14'd 16373;
        11'd 24:out = 14'd 16372;
        11'd 25:out = 14'd 16371;
        11'd 26:out = 14'd 16370;
        11'd 27:out = 14'd 16369;
        11'd 28:out = 14'd 16368;
        11'd 29:out = 14'd 16367;
        11'd 30:out = 14'd 16366;
        11'd 31:out = 14'd 16365;
        11'd 32:out = 14'd 16364;
        11'd 33:out = 14'd 16363;
        11'd 34:out = 14'd 16361;
        11'd 35:out = 14'd 16360;
        11'd 36:out = 14'd 16359;
        11'd 37:out = 14'd 16357;
        11'd 38:out = 14'd 16356;
        11'd 39:out = 14'd 16354;
        11'd 40:out = 14'd 16353;
        11'd 41:out = 14'd 16351;
        11'd 42:out = 14'd 16350;
        11'd 43:out = 14'd 16348;
        11'd 44:out = 14'd 16346;
        11'd 45:out = 14'd 16344;
        11'd 46:out = 14'd 16343;
        11'd 47:out = 14'd 16341;
        11'd 48:out = 14'd 16339;
        11'd 49:out = 14'd 16337;
        11'd 50:out = 14'd 16335;
        11'd 51:out = 14'd 16333;
        11'd 52:out = 14'd 16331;
        11'd 53:out = 14'd 16329;
        11'd 54:out = 14'd 16327;
        11'd 55:out = 14'd 16325;
        11'd 56:out = 14'd 16323;
        11'd 57:out = 14'd 16321;
        11'd 58:out = 14'd 16319;
        11'd 59:out = 14'd 16316;
        11'd 60:out = 14'd 16314;
        11'd 61:out = 14'd 16312;
        11'd 62:out = 14'd 16309;
        11'd 63:out = 14'd 16307;
        11'd 64:out = 14'd 16305;
        11'd 65:out = 14'd 16302;
        11'd 66:out = 14'd 16300;
        11'd 67:out = 14'd 16297;
        11'd 68:out = 14'd 16294;
        11'd 69:out = 14'd 16292;
        11'd 70:out = 14'd 16289;
        11'd 71:out = 14'd 16286;
        11'd 72:out = 14'd 16284;
        11'd 73:out = 14'd 16281;
        11'd 74:out = 14'd 16278;
        11'd 75:out = 14'd 16275;
        11'd 76:out = 14'd 16272;
        11'd 77:out = 14'd 16269;
        11'd 78:out = 14'd 16266;
        11'd 79:out = 14'd 16263;
        11'd 80:out = 14'd 16260;
        11'd 81:out = 14'd 16257;
        11'd 82:out = 14'd 16254;
        11'd 83:out = 14'd 16251;
        11'd 84:out = 14'd 16248;
        11'd 85:out = 14'd 16244;
        11'd 86:out = 14'd 16241;
        11'd 87:out = 14'd 16238;
        11'd 88:out = 14'd 16234;
        11'd 89:out = 14'd 16231;
        11'd 90:out = 14'd 16228;
        11'd 91:out = 14'd 16224;
        11'd 92:out = 14'd 16221;
        11'd 93:out = 14'd 16217;
        11'd 94:out = 14'd 16213;
        11'd 95:out = 14'd 16210;
        11'd 96:out = 14'd 16206;
        11'd 97:out = 14'd 16202;
        11'd 98:out = 14'd 16199;
        11'd 99:out = 14'd 16195;
        11'd 100:out = 14'd 16191;
        11'd 101:out = 14'd 16187;
        11'd 102:out = 14'd 16183;
        11'd 103:out = 14'd 16179;
        11'd 104:out = 14'd 16175;
        11'd 105:out = 14'd 16171;
        11'd 106:out = 14'd 16167;
        11'd 107:out = 14'd 16163;
        11'd 108:out = 14'd 16159;
        11'd 109:out = 14'd 16155;
        11'd 110:out = 14'd 16151;
        11'd 111:out = 14'd 16147;
        11'd 112:out = 14'd 16142;
        11'd 113:out = 14'd 16138;
        11'd 114:out = 14'd 16134;
        11'd 115:out = 14'd 16129;
        11'd 116:out = 14'd 16125;
        11'd 117:out = 14'd 16120;
        11'd 118:out = 14'd 16116;
        11'd 119:out = 14'd 16111;
        11'd 120:out = 14'd 16107;
        11'd 121:out = 14'd 16102;
        11'd 122:out = 14'd 16097;
        11'd 123:out = 14'd 16093;
        11'd 124:out = 14'd 16088;
        11'd 125:out = 14'd 16083;
        11'd 126:out = 14'd 16078;
        11'd 127:out = 14'd 16074;
        11'd 128:out = 14'd 16069;
        11'd 129:out = 14'd 16064;
        11'd 130:out = 14'd 16059;
        11'd 131:out = 14'd 16054;
        11'd 132:out = 14'd 16049;
        11'd 133:out = 14'd 16044;
        11'd 134:out = 14'd 16039;
        11'd 135:out = 14'd 16033;
        11'd 136:out = 14'd 16028;
        11'd 137:out = 14'd 16023;
        11'd 138:out = 14'd 16018;
        11'd 139:out = 14'd 16012;
        11'd 140:out = 14'd 16007;
        11'd 141:out = 14'd 16002;
        11'd 142:out = 14'd 15996;
        11'd 143:out = 14'd 15991;
        11'd 144:out = 14'd 15985;
        11'd 145:out = 14'd 15980;
        11'd 146:out = 14'd 15974;
        11'd 147:out = 14'd 15969;
        11'd 148:out = 14'd 15963;
        11'd 149:out = 14'd 15957;
        11'd 150:out = 14'd 15952;
        11'd 151:out = 14'd 15946;
        11'd 152:out = 14'd 15940;
        11'd 153:out = 14'd 15934;
        11'd 154:out = 14'd 15928;
        11'd 155:out = 14'd 15923;
        11'd 156:out = 14'd 15917;
        11'd 157:out = 14'd 15911;
        11'd 158:out = 14'd 15905;
        11'd 159:out = 14'd 15899;
        11'd 160:out = 14'd 15892;
        11'd 161:out = 14'd 15886;
        11'd 162:out = 14'd 15880;
        11'd 163:out = 14'd 15874;
        11'd 164:out = 14'd 15868;
        11'd 165:out = 14'd 15861;
        11'd 166:out = 14'd 15855;
        11'd 167:out = 14'd 15849;
        11'd 168:out = 14'd 15842;
        11'd 169:out = 14'd 15836;
        11'd 170:out = 14'd 15830;
        11'd 171:out = 14'd 15823;
        11'd 172:out = 14'd 15817;
        11'd 173:out = 14'd 15810;
        11'd 174:out = 14'd 15803;
        11'd 175:out = 14'd 15797;
        11'd 176:out = 14'd 15790;
        11'd 177:out = 14'd 15783;
        11'd 178:out = 14'd 15777;
        11'd 179:out = 14'd 15770;
        11'd 180:out = 14'd 15763;
        11'd 181:out = 14'd 15756;
        11'd 182:out = 14'd 15749;
        11'd 183:out = 14'd 15742;
        11'd 184:out = 14'd 15735;
        11'd 185:out = 14'd 15728;
        11'd 186:out = 14'd 15721;
        11'd 187:out = 14'd 15714;
        11'd 188:out = 14'd 15707;
        11'd 189:out = 14'd 15700;
        11'd 190:out = 14'd 15693;
        11'd 191:out = 14'd 15685;
        11'd 192:out = 14'd 15678;
        11'd 193:out = 14'd 15671;
        11'd 194:out = 14'd 15663;
        11'd 195:out = 14'd 15656;
        11'd 196:out = 14'd 15649;
        11'd 197:out = 14'd 15641;
        11'd 198:out = 14'd 15634;
        11'd 199:out = 14'd 15626;
        11'd 200:out = 14'd 15618;
        11'd 201:out = 14'd 15611;
        11'd 202:out = 14'd 15603;
        11'd 203:out = 14'd 15596;
        11'd 204:out = 14'd 15588;
        11'd 205:out = 14'd 15580;
        11'd 206:out = 14'd 15572;
        11'd 207:out = 14'd 15564;
        11'd 208:out = 14'd 15557;
        11'd 209:out = 14'd 15549;
        11'd 210:out = 14'd 15541;
        11'd 211:out = 14'd 15533;
        11'd 212:out = 14'd 15525;
        11'd 213:out = 14'd 15517;
        11'd 214:out = 14'd 15509;
        11'd 215:out = 14'd 15500;
        11'd 216:out = 14'd 15492;
        11'd 217:out = 14'd 15484;
        11'd 218:out = 14'd 15476;
        11'd 219:out = 14'd 15468;
        11'd 220:out = 14'd 15459;
        11'd 221:out = 14'd 15451;
        11'd 222:out = 14'd 15443;
        11'd 223:out = 14'd 15434;
        11'd 224:out = 14'd 15426;
        11'd 225:out = 14'd 15417;
        11'd 226:out = 14'd 15409;
        11'd 227:out = 14'd 15400;
        11'd 228:out = 14'd 15392;
        11'd 229:out = 14'd 15383;
        11'd 230:out = 14'd 15374;
        11'd 231:out = 14'd 15366;
        11'd 232:out = 14'd 15357;
        11'd 233:out = 14'd 15348;
        11'd 234:out = 14'd 15339;
        11'd 235:out = 14'd 15330;
        11'd 236:out = 14'd 15322;
        11'd 237:out = 14'd 15313;
        11'd 238:out = 14'd 15304;
        11'd 239:out = 14'd 15295;
        11'd 240:out = 14'd 15286;
        11'd 241:out = 14'd 15277;
        11'd 242:out = 14'd 15267;
        11'd 243:out = 14'd 15258;
        11'd 244:out = 14'd 15249;
        11'd 245:out = 14'd 15240;
        11'd 246:out = 14'd 15231;
        11'd 247:out = 14'd 15221;
        11'd 248:out = 14'd 15212;
        11'd 249:out = 14'd 15203;
        11'd 250:out = 14'd 15193;
        11'd 251:out = 14'd 15184;
        11'd 252:out = 14'd 15175;
        11'd 253:out = 14'd 15165;
        11'd 254:out = 14'd 15156;
        11'd 255:out = 14'd 15146;
        11'd 256:out = 14'd 15136;
        11'd 257:out = 14'd 15127;
        11'd 258:out = 14'd 15117;
        11'd 259:out = 14'd 15107;
        11'd 260:out = 14'd 15098;
        11'd 261:out = 14'd 15088;
        11'd 262:out = 14'd 15078;
        11'd 263:out = 14'd 15068;
        11'd 264:out = 14'd 15058;
        11'd 265:out = 14'd 15048;
        11'd 266:out = 14'd 15038;
        11'd 267:out = 14'd 15028;
        11'd 268:out = 14'd 15018;
        11'd 269:out = 14'd 15008;
        11'd 270:out = 14'd 14998;
        11'd 271:out = 14'd 14988;
        11'd 272:out = 14'd 14978;
        11'd 273:out = 14'd 14968;
        11'd 274:out = 14'd 14957;
        11'd 275:out = 14'd 14947;
        11'd 276:out = 14'd 14937;
        11'd 277:out = 14'd 14927;
        11'd 278:out = 14'd 14916;
        11'd 279:out = 14'd 14906;
        11'd 280:out = 14'd 14895;
        11'd 281:out = 14'd 14885;
        11'd 282:out = 14'd 14874;
        11'd 283:out = 14'd 14864;
        11'd 284:out = 14'd 14853;
        11'd 285:out = 14'd 14843;
        11'd 286:out = 14'd 14832;
        11'd 287:out = 14'd 14821;
        11'd 288:out = 14'd 14810;
        11'd 289:out = 14'd 14800;
        11'd 290:out = 14'd 14789;
        11'd 291:out = 14'd 14778;
        11'd 292:out = 14'd 14767;
        11'd 293:out = 14'd 14756;
        11'd 294:out = 14'd 14745;
        11'd 295:out = 14'd 14734;
        11'd 296:out = 14'd 14723;
        11'd 297:out = 14'd 14712;
        11'd 298:out = 14'd 14701;
        11'd 299:out = 14'd 14690;
        11'd 300:out = 14'd 14679;
        11'd 301:out = 14'd 14668;
        11'd 302:out = 14'd 14657;
        11'd 303:out = 14'd 14645;
        11'd 304:out = 14'd 14634;
        11'd 305:out = 14'd 14623;
        11'd 306:out = 14'd 14611;
        11'd 307:out = 14'd 14600;
        11'd 308:out = 14'd 14589;
        11'd 309:out = 14'd 14577;
        11'd 310:out = 14'd 14566;
        11'd 311:out = 14'd 14554;
        11'd 312:out = 14'd 14543;
        11'd 313:out = 14'd 14531;
        11'd 314:out = 14'd 14519;
        11'd 315:out = 14'd 14508;
        11'd 316:out = 14'd 14496;
        11'd 317:out = 14'd 14484;
        11'd 318:out = 14'd 14473;
        11'd 319:out = 14'd 14461;
        11'd 320:out = 14'd 14449;
        11'd 321:out = 14'd 14437;
        11'd 322:out = 14'd 14425;
        11'd 323:out = 14'd 14413;
        11'd 324:out = 14'd 14401;
        11'd 325:out = 14'd 14389;
        11'd 326:out = 14'd 14377;
        11'd 327:out = 14'd 14365;
        11'd 328:out = 14'd 14353;
        11'd 329:out = 14'd 14341;
        11'd 330:out = 14'd 14329;
        11'd 331:out = 14'd 14317;
        11'd 332:out = 14'd 14304;
        11'd 333:out = 14'd 14292;
        11'd 334:out = 14'd 14280;
        11'd 335:out = 14'd 14267;
        11'd 336:out = 14'd 14255;
        11'd 337:out = 14'd 14243;
        11'd 338:out = 14'd 14230;
        11'd 339:out = 14'd 14218;
        11'd 340:out = 14'd 14205;
        11'd 341:out = 14'd 14193;
        11'd 342:out = 14'd 14180;
        11'd 343:out = 14'd 14167;
        11'd 344:out = 14'd 14155;
        11'd 345:out = 14'd 14142;
        11'd 346:out = 14'd 14129;
        11'd 347:out = 14'd 14117;
        11'd 348:out = 14'd 14104;
        11'd 349:out = 14'd 14091;
        11'd 350:out = 14'd 14078;
        11'd 351:out = 14'd 14065;
        11'd 352:out = 14'd 14053;
        11'd 353:out = 14'd 14040;
        11'd 354:out = 14'd 14027;
        11'd 355:out = 14'd 14014;
        11'd 356:out = 14'd 14001;
        11'd 357:out = 14'd 13988;
        11'd 358:out = 14'd 13974;
        11'd 359:out = 14'd 13961;
        11'd 360:out = 14'd 13948;
        11'd 361:out = 14'd 13935;
        11'd 362:out = 14'd 13922;
        11'd 363:out = 14'd 13908;
        11'd 364:out = 14'd 13895;
        11'd 365:out = 14'd 13882;
        11'd 366:out = 14'd 13868;
        11'd 367:out = 14'd 13855;
        11'd 368:out = 14'd 13842;
        11'd 369:out = 14'd 13828;
        11'd 370:out = 14'd 13815;
        11'd 371:out = 14'd 13801;
        11'd 372:out = 14'd 13788;
        11'd 373:out = 14'd 13774;
        11'd 374:out = 14'd 13760;
        11'd 375:out = 14'd 13747;
        11'd 376:out = 14'd 13733;
        11'd 377:out = 14'd 13719;
        11'd 378:out = 14'd 13705;
        11'd 379:out = 14'd 13692;
        11'd 380:out = 14'd 13678;
        11'd 381:out = 14'd 13664;
        11'd 382:out = 14'd 13650;
        11'd 383:out = 14'd 13636;
        11'd 384:out = 14'd 13622;
        11'd 385:out = 14'd 13608;
        11'd 386:out = 14'd 13594;
        11'd 387:out = 14'd 13580;
        11'd 388:out = 14'd 13566;
        11'd 389:out = 14'd 13552;
        11'd 390:out = 14'd 13538;
        11'd 391:out = 14'd 13524;
        11'd 392:out = 14'd 13510;
        11'd 393:out = 14'd 13495;
        11'd 394:out = 14'd 13481;
        11'd 395:out = 14'd 13467;
        11'd 396:out = 14'd 13452;
        11'd 397:out = 14'd 13438;
        11'd 398:out = 14'd 13424;
        11'd 399:out = 14'd 13409;
        11'd 400:out = 14'd 13395;
        11'd 401:out = 14'd 13380;
        11'd 402:out = 14'd 13366;
        11'd 403:out = 14'd 13351;
        11'd 404:out = 14'd 13337;
        11'd 405:out = 14'd 13322;
        11'd 406:out = 14'd 13307;
        11'd 407:out = 14'd 13293;
        11'd 408:out = 14'd 13278;
        11'd 409:out = 14'd 13263;
        11'd 410:out = 14'd 13249;
        11'd 411:out = 14'd 13234;
        11'd 412:out = 14'd 13219;
        11'd 413:out = 14'd 13204;
        11'd 414:out = 14'd 13189;
        11'd 415:out = 14'd 13174;
        11'd 416:out = 14'd 13159;
        11'd 417:out = 14'd 13144;
        11'd 418:out = 14'd 13129;
        11'd 419:out = 14'd 13114;
        11'd 420:out = 14'd 13099;
        11'd 421:out = 14'd 13084;
        11'd 422:out = 14'd 13069;
        11'd 423:out = 14'd 13054;
        11'd 424:out = 14'd 13038;
        11'd 425:out = 14'd 13023;
        11'd 426:out = 14'd 13008;
        11'd 427:out = 14'd 12993;
        11'd 428:out = 14'd 12977;
        11'd 429:out = 14'd 12962;
        11'd 430:out = 14'd 12947;
        11'd 431:out = 14'd 12931;
        11'd 432:out = 14'd 12916;
        11'd 433:out = 14'd 12900;
        11'd 434:out = 14'd 12885;
        11'd 435:out = 14'd 12869;
        11'd 436:out = 14'd 12854;
        11'd 437:out = 14'd 12838;
        11'd 438:out = 14'd 12822;
        11'd 439:out = 14'd 12807;
        11'd 440:out = 14'd 12791;
        11'd 441:out = 14'd 12775;
        11'd 442:out = 14'd 12760;
        11'd 443:out = 14'd 12744;
        11'd 444:out = 14'd 12728;
        11'd 445:out = 14'd 12712;
        11'd 446:out = 14'd 12696;
        11'd 447:out = 14'd 12680;
        11'd 448:out = 14'd 12665;
        11'd 449:out = 14'd 12649;
        11'd 450:out = 14'd 12633;
        11'd 451:out = 14'd 12617;
        11'd 452:out = 14'd 12600;
        11'd 453:out = 14'd 12584;
        11'd 454:out = 14'd 12568;
        11'd 455:out = 14'd 12552;
        11'd 456:out = 14'd 12536;
        11'd 457:out = 14'd 12520;
        11'd 458:out = 14'd 12504;
        11'd 459:out = 14'd 12487;
        11'd 460:out = 14'd 12471;
        11'd 461:out = 14'd 12455;
        11'd 462:out = 14'd 12438;
        11'd 463:out = 14'd 12422;
        11'd 464:out = 14'd 12406;
        11'd 465:out = 14'd 12389;
        11'd 466:out = 14'd 12373;
        11'd 467:out = 14'd 12356;
        11'd 468:out = 14'd 12340;
        11'd 469:out = 14'd 12323;
        11'd 470:out = 14'd 12307;
        11'd 471:out = 14'd 12290;
        11'd 472:out = 14'd 12273;
        11'd 473:out = 14'd 12257;
        11'd 474:out = 14'd 12240;
        11'd 475:out = 14'd 12223;
        11'd 476:out = 14'd 12207;
        11'd 477:out = 14'd 12190;
        11'd 478:out = 14'd 12173;
        11'd 479:out = 14'd 12156;
        11'd 480:out = 14'd 12139;
        11'd 481:out = 14'd 12122;
        11'd 482:out = 14'd 12105;
        11'd 483:out = 14'd 12088;
        11'd 484:out = 14'd 12072;
        11'd 485:out = 14'd 12054;
        11'd 486:out = 14'd 12037;
        11'd 487:out = 14'd 12020;
        11'd 488:out = 14'd 12003;
        11'd 489:out = 14'd 11986;
        11'd 490:out = 14'd 11969;
        11'd 491:out = 14'd 11952;
        11'd 492:out = 14'd 11935;
        11'd 493:out = 14'd 11917;
        11'd 494:out = 14'd 11900;
        11'd 495:out = 14'd 11883;
        11'd 496:out = 14'd 11866;
        11'd 497:out = 14'd 11848;
        11'd 498:out = 14'd 11831;
        11'd 499:out = 14'd 11813;
        11'd 500:out = 14'd 11796;
        11'd 501:out = 14'd 11779;
        11'd 502:out = 14'd 11761;
        11'd 503:out = 14'd 11744;
        11'd 504:out = 14'd 11726;
        11'd 505:out = 14'd 11708;
        11'd 506:out = 14'd 11691;
        11'd 507:out = 14'd 11673;
        11'd 508:out = 14'd 11656;
        11'd 509:out = 14'd 11638;
        11'd 510:out = 14'd 11620;
        11'd 511:out = 14'd 11602;
        11'd 512:out = 14'd 11585;
        11'd 513:out = 14'd 11567;
        11'd 514:out = 14'd 11549;
        11'd 515:out = 14'd 11531;
        11'd 516:out = 14'd 11513;
        11'd 517:out = 14'd 11496;
        11'd 518:out = 14'd 11478;
        11'd 519:out = 14'd 11460;
        11'd 520:out = 14'd 11442;
        11'd 521:out = 14'd 11424;
        11'd 522:out = 14'd 11406;
        11'd 523:out = 14'd 11388;
        11'd 524:out = 14'd 11370;
        11'd 525:out = 14'd 11351;
        11'd 526:out = 14'd 11333;
        11'd 527:out = 14'd 11315;
        11'd 528:out = 14'd 11297;
        11'd 529:out = 14'd 11279;
        11'd 530:out = 14'd 11260;
        11'd 531:out = 14'd 11242;
        11'd 532:out = 14'd 11224;
        11'd 533:out = 14'd 11206;
        11'd 534:out = 14'd 11187;
        11'd 535:out = 14'd 11169;
        11'd 536:out = 14'd 11150;
        11'd 537:out = 14'd 11132;
        11'd 538:out = 14'd 11114;
        11'd 539:out = 14'd 11095;
        11'd 540:out = 14'd 11077;
        11'd 541:out = 14'd 11058;
        11'd 542:out = 14'd 11040;
        11'd 543:out = 14'd 11021;
        11'd 544:out = 14'd 11002;
        11'd 545:out = 14'd 10984;
        11'd 546:out = 14'd 10965;
        11'd 547:out = 14'd 10946;
        11'd 548:out = 14'd 10928;
        11'd 549:out = 14'd 10909;
        11'd 550:out = 14'd 10890;
        11'd 551:out = 14'd 10871;
        11'd 552:out = 14'd 10853;
        11'd 553:out = 14'd 10834;
        11'd 554:out = 14'd 10815;
        11'd 555:out = 14'd 10796;
        11'd 556:out = 14'd 10777;
        11'd 557:out = 14'd 10758;
        11'd 558:out = 14'd 10739;
        11'd 559:out = 14'd 10720;
        11'd 560:out = 14'd 10701;
        11'd 561:out = 14'd 10682;
        11'd 562:out = 14'd 10663;
        11'd 563:out = 14'd 10644;
        11'd 564:out = 14'd 10625;
        11'd 565:out = 14'd 10606;
        11'd 566:out = 14'd 10586;
        11'd 567:out = 14'd 10567;
        11'd 568:out = 14'd 10548;
        11'd 569:out = 14'd 10529;
        11'd 570:out = 14'd 10510;
        11'd 571:out = 14'd 10490;
        11'd 572:out = 14'd 10471;
        11'd 573:out = 14'd 10452;
        11'd 574:out = 14'd 10432;
        11'd 575:out = 14'd 10413;
        11'd 576:out = 14'd 10393;
        11'd 577:out = 14'd 10374;
        11'd 578:out = 14'd 10354;
        11'd 579:out = 14'd 10335;
        11'd 580:out = 14'd 10315;
        11'd 581:out = 14'd 10296;
        11'd 582:out = 14'd 10276;
        11'd 583:out = 14'd 10257;
        11'd 584:out = 14'd 10237;
        11'd 585:out = 14'd 10218;
        11'd 586:out = 14'd 10198;
        11'd 587:out = 14'd 10178;
        11'd 588:out = 14'd 10159;
        11'd 589:out = 14'd 10139;
        11'd 590:out = 14'd 10119;
        11'd 591:out = 14'd 10099;
        11'd 592:out = 14'd 10079;
        11'd 593:out = 14'd 10060;
        11'd 594:out = 14'd 10040;
        11'd 595:out = 14'd 10020;
        11'd 596:out = 14'd 10000;
        11'd 597:out = 14'd 9980;
        11'd 598:out = 14'd 9960;
        11'd 599:out = 14'd 9940;
        11'd 600:out = 14'd 9920;
        11'd 601:out = 14'd 9900;
        11'd 602:out = 14'd 9880;
        11'd 603:out = 14'd 9860;
        11'd 604:out = 14'd 9840;
        11'd 605:out = 14'd 9820;
        11'd 606:out = 14'd 9800;
        11'd 607:out = 14'd 9780;
        11'd 608:out = 14'd 9759;
        11'd 609:out = 14'd 9739;
        11'd 610:out = 14'd 9719;
        11'd 611:out = 14'd 9699;
        11'd 612:out = 14'd 9679;
        11'd 613:out = 14'd 9658;
        11'd 614:out = 14'd 9638;
        11'd 615:out = 14'd 9618;
        11'd 616:out = 14'd 9597;
        11'd 617:out = 14'd 9577;
        11'd 618:out = 14'd 9556;
        11'd 619:out = 14'd 9536;
        11'd 620:out = 14'd 9516;
        11'd 621:out = 14'd 9495;
        11'd 622:out = 14'd 9475;
        11'd 623:out = 14'd 9454;
        11'd 624:out = 14'd 9434;
        11'd 625:out = 14'd 9413;
        11'd 626:out = 14'd 9392;
        11'd 627:out = 14'd 9372;
        11'd 628:out = 14'd 9351;
        11'd 629:out = 14'd 9331;
        11'd 630:out = 14'd 9310;
        11'd 631:out = 14'd 9289;
        11'd 632:out = 14'd 9268;
        11'd 633:out = 14'd 9248;
        11'd 634:out = 14'd 9227;
        11'd 635:out = 14'd 9206;
        11'd 636:out = 14'd 9185;
        11'd 637:out = 14'd 9165;
        11'd 638:out = 14'd 9144;
        11'd 639:out = 14'd 9123;
        11'd 640:out = 14'd 9102;
        11'd 641:out = 14'd 9081;
        11'd 642:out = 14'd 9060;
        11'd 643:out = 14'd 9039;
        11'd 644:out = 14'd 9018;
        11'd 645:out = 14'd 8997;
        11'd 646:out = 14'd 8976;
        11'd 647:out = 14'd 8955;
        11'd 648:out = 14'd 8934;
        11'd 649:out = 14'd 8913;
        11'd 650:out = 14'd 8892;
        11'd 651:out = 14'd 8871;
        11'd 652:out = 14'd 8850;
        11'd 653:out = 14'd 8829;
        11'd 654:out = 14'd 8807;
        11'd 655:out = 14'd 8786;
        11'd 656:out = 14'd 8765;
        11'd 657:out = 14'd 8744;
        11'd 658:out = 14'd 8722;
        11'd 659:out = 14'd 8701;
        11'd 660:out = 14'd 8680;
        11'd 661:out = 14'd 8658;
        11'd 662:out = 14'd 8637;
        11'd 663:out = 14'd 8616;
        11'd 664:out = 14'd 8594;
        11'd 665:out = 14'd 8573;
        11'd 666:out = 14'd 8552;
        11'd 667:out = 14'd 8530;
        11'd 668:out = 14'd 8509;
        11'd 669:out = 14'd 8487;
        11'd 670:out = 14'd 8466;
        11'd 671:out = 14'd 8444;
        11'd 672:out = 14'd 8423;
        11'd 673:out = 14'd 8401;
        11'd 674:out = 14'd 8379;
        11'd 675:out = 14'd 8358;
        11'd 676:out = 14'd 8336;
        11'd 677:out = 14'd 8315;
        11'd 678:out = 14'd 8293;
        11'd 679:out = 14'd 8271;
        11'd 680:out = 14'd 8249;
        11'd 681:out = 14'd 8228;
        11'd 682:out = 14'd 8206;
        11'd 683:out = 14'd 8184;
        11'd 684:out = 14'd 8162;
        11'd 685:out = 14'd 8141;
        11'd 686:out = 14'd 8119;
        11'd 687:out = 14'd 8097;
        11'd 688:out = 14'd 8075;
        11'd 689:out = 14'd 8053;
        11'd 690:out = 14'd 8031;
        11'd 691:out = 14'd 8009;
        11'd 692:out = 14'd 7988;
        11'd 693:out = 14'd 7966;
        11'd 694:out = 14'd 7944;
        11'd 695:out = 14'd 7922;
        11'd 696:out = 14'd 7900;
        11'd 697:out = 14'd 7878;
        11'd 698:out = 14'd 7856;
        11'd 699:out = 14'd 7833;
        11'd 700:out = 14'd 7811;
        11'd 701:out = 14'd 7789;
        11'd 702:out = 14'd 7767;
        11'd 703:out = 14'd 7745;
        11'd 704:out = 14'd 7723;
        11'd 705:out = 14'd 7701;
        11'd 706:out = 14'd 7678;
        11'd 707:out = 14'd 7656;
        11'd 708:out = 14'd 7634;
        11'd 709:out = 14'd 7612;
        11'd 710:out = 14'd 7590;
        11'd 711:out = 14'd 7567;
        11'd 712:out = 14'd 7545;
        11'd 713:out = 14'd 7523;
        11'd 714:out = 14'd 7500;
        11'd 715:out = 14'd 7478;
        11'd 716:out = 14'd 7456;
        11'd 717:out = 14'd 7433;
        11'd 718:out = 14'd 7411;
        11'd 719:out = 14'd 7388;
        11'd 720:out = 14'd 7366;
        11'd 721:out = 14'd 7343;
        11'd 722:out = 14'd 7321;
        11'd 723:out = 14'd 7299;
        11'd 724:out = 14'd 7276;
        11'd 725:out = 14'd 7253;
        11'd 726:out = 14'd 7231;
        11'd 727:out = 14'd 7208;
        11'd 728:out = 14'd 7186;
        11'd 729:out = 14'd 7163;
        11'd 730:out = 14'd 7141;
        11'd 731:out = 14'd 7118;
        11'd 732:out = 14'd 7095;
        11'd 733:out = 14'd 7073;
        11'd 734:out = 14'd 7050;
        11'd 735:out = 14'd 7027;
        11'd 736:out = 14'd 7005;
        11'd 737:out = 14'd 6982;
        11'd 738:out = 14'd 6959;
        11'd 739:out = 14'd 6936;
        11'd 740:out = 14'd 6914;
        11'd 741:out = 14'd 6891;
        11'd 742:out = 14'd 6868;
        11'd 743:out = 14'd 6845;
        11'd 744:out = 14'd 6822;
        11'd 745:out = 14'd 6799;
        11'd 746:out = 14'd 6777;
        11'd 747:out = 14'd 6754;
        11'd 748:out = 14'd 6731;
        11'd 749:out = 14'd 6708;
        11'd 750:out = 14'd 6685;
        11'd 751:out = 14'd 6662;
        11'd 752:out = 14'd 6639;
        11'd 753:out = 14'd 6616;
        11'd 754:out = 14'd 6593;
        11'd 755:out = 14'd 6570;
        11'd 756:out = 14'd 6547;
        11'd 757:out = 14'd 6524;
        11'd 758:out = 14'd 6501;
        11'd 759:out = 14'd 6478;
        11'd 760:out = 14'd 6455;
        11'd 761:out = 14'd 6432;
        11'd 762:out = 14'd 6408;
        11'd 763:out = 14'd 6385;
        11'd 764:out = 14'd 6362;
        11'd 765:out = 14'd 6339;
        11'd 766:out = 14'd 6316;
        11'd 767:out = 14'd 6293;
        11'd 768:out = 14'd 6269;
        11'd 769:out = 14'd 6246;
        11'd 770:out = 14'd 6223;
        11'd 771:out = 14'd 6200;
        11'd 772:out = 14'd 6176;
        11'd 773:out = 14'd 6153;
        11'd 774:out = 14'd 6130;
        11'd 775:out = 14'd 6106;
        11'd 776:out = 14'd 6083;
        11'd 777:out = 14'd 6060;
        11'd 778:out = 14'd 6036;
        11'd 779:out = 14'd 6013;
        11'd 780:out = 14'd 5990;
        11'd 781:out = 14'd 5966;
        11'd 782:out = 14'd 5943;
        11'd 783:out = 14'd 5919;
        11'd 784:out = 14'd 5896;
        11'd 785:out = 14'd 5873;
        11'd 786:out = 14'd 5849;
        11'd 787:out = 14'd 5826;
        11'd 788:out = 14'd 5802;
        11'd 789:out = 14'd 5779;
        11'd 790:out = 14'd 5755;
        11'd 791:out = 14'd 5732;
        11'd 792:out = 14'd 5708;
        11'd 793:out = 14'd 5684;
        11'd 794:out = 14'd 5661;
        11'd 795:out = 14'd 5637;
        11'd 796:out = 14'd 5614;
        11'd 797:out = 14'd 5590;
        11'd 798:out = 14'd 5566;
        11'd 799:out = 14'd 5543;
        11'd 800:out = 14'd 5519;
        11'd 801:out = 14'd 5495;
        11'd 802:out = 14'd 5472;
        11'd 803:out = 14'd 5448;
        11'd 804:out = 14'd 5424;
        11'd 805:out = 14'd 5401;
        11'd 806:out = 14'd 5377;
        11'd 807:out = 14'd 5353;
        11'd 808:out = 14'd 5329;
        11'd 809:out = 14'd 5306;
        11'd 810:out = 14'd 5282;
        11'd 811:out = 14'd 5258;
        11'd 812:out = 14'd 5234;
        11'd 813:out = 14'd 5210;
        11'd 814:out = 14'd 5187;
        11'd 815:out = 14'd 5163;
        11'd 816:out = 14'd 5139;
        11'd 817:out = 14'd 5115;
        11'd 818:out = 14'd 5091;
        11'd 819:out = 14'd 5067;
        11'd 820:out = 14'd 5043;
        11'd 821:out = 14'd 5019;
        11'd 822:out = 14'd 4995;
        11'd 823:out = 14'd 4972;
        11'd 824:out = 14'd 4948;
        11'd 825:out = 14'd 4924;
        11'd 826:out = 14'd 4900;
        11'd 827:out = 14'd 4876;
        11'd 828:out = 14'd 4852;
        11'd 829:out = 14'd 4828;
        11'd 830:out = 14'd 4804;
        11'd 831:out = 14'd 4780;
        11'd 832:out = 14'd 4756;
        11'd 833:out = 14'd 4731;
        11'd 834:out = 14'd 4707;
        11'd 835:out = 14'd 4683;
        11'd 836:out = 14'd 4659;
        11'd 837:out = 14'd 4635;
        11'd 838:out = 14'd 4611;
        11'd 839:out = 14'd 4587;
        11'd 840:out = 14'd 4563;
        11'd 841:out = 14'd 4539;
        11'd 842:out = 14'd 4514;
        11'd 843:out = 14'd 4490;
        11'd 844:out = 14'd 4466;
        11'd 845:out = 14'd 4442;
        11'd 846:out = 14'd 4418;
        11'd 847:out = 14'd 4394;
        11'd 848:out = 14'd 4369;
        11'd 849:out = 14'd 4345;
        11'd 850:out = 14'd 4321;
        11'd 851:out = 14'd 4297;
        11'd 852:out = 14'd 4272;
        11'd 853:out = 14'd 4248;
        11'd 854:out = 14'd 4224;
        11'd 855:out = 14'd 4200;
        11'd 856:out = 14'd 4175;
        11'd 857:out = 14'd 4151;
        11'd 858:out = 14'd 4127;
        11'd 859:out = 14'd 4102;
        11'd 860:out = 14'd 4078;
        11'd 861:out = 14'd 4054;
        11'd 862:out = 14'd 4029;
        11'd 863:out = 14'd 4005;
        11'd 864:out = 14'd 3980;
        11'd 865:out = 14'd 3956;
        11'd 866:out = 14'd 3932;
        11'd 867:out = 14'd 3907;
        11'd 868:out = 14'd 3883;
        11'd 869:out = 14'd 3858;
        11'd 870:out = 14'd 3834;
        11'd 871:out = 14'd 3810;
        11'd 872:out = 14'd 3785;
        11'd 873:out = 14'd 3761;
        11'd 874:out = 14'd 3736;
        11'd 875:out = 14'd 3712;
        11'd 876:out = 14'd 3687;
        11'd 877:out = 14'd 3663;
        11'd 878:out = 14'd 3638;
        11'd 879:out = 14'd 3614;
        11'd 880:out = 14'd 3589;
        11'd 881:out = 14'd 3565;
        11'd 882:out = 14'd 3540;
        11'd 883:out = 14'd 3516;
        11'd 884:out = 14'd 3491;
        11'd 885:out = 14'd 3467;
        11'd 886:out = 14'd 3442;
        11'd 887:out = 14'd 3417;
        11'd 888:out = 14'd 3393;
        11'd 889:out = 14'd 3368;
        11'd 890:out = 14'd 3344;
        11'd 891:out = 14'd 3319;
        11'd 892:out = 14'd 3294;
        11'd 893:out = 14'd 3270;
        11'd 894:out = 14'd 3245;
        11'd 895:out = 14'd 3221;
        11'd 896:out = 14'd 3196;
        11'd 897:out = 14'd 3171;
        11'd 898:out = 14'd 3147;
        11'd 899:out = 14'd 3122;
        11'd 900:out = 14'd 3097;
        11'd 901:out = 14'd 3073;
        11'd 902:out = 14'd 3048;
        11'd 903:out = 14'd 3023;
        11'd 904:out = 14'd 2998;
        11'd 905:out = 14'd 2974;
        11'd 906:out = 14'd 2949;
        11'd 907:out = 14'd 2924;
        11'd 908:out = 14'd 2900;
        11'd 909:out = 14'd 2875;
        11'd 910:out = 14'd 2850;
        11'd 911:out = 14'd 2825;
        11'd 912:out = 14'd 2801;
        11'd 913:out = 14'd 2776;
        11'd 914:out = 14'd 2751;
        11'd 915:out = 14'd 2726;
        11'd 916:out = 14'd 2701;
        11'd 917:out = 14'd 2677;
        11'd 918:out = 14'd 2652;
        11'd 919:out = 14'd 2627;
        11'd 920:out = 14'd 2602;
        11'd 921:out = 14'd 2577;
        11'd 922:out = 14'd 2553;
        11'd 923:out = 14'd 2528;
        11'd 924:out = 14'd 2503;
        11'd 925:out = 14'd 2478;
        11'd 926:out = 14'd 2453;
        11'd 927:out = 14'd 2428;
        11'd 928:out = 14'd 2404;
        11'd 929:out = 14'd 2379;
        11'd 930:out = 14'd 2354;
        11'd 931:out = 14'd 2329;
        11'd 932:out = 14'd 2304;
        11'd 933:out = 14'd 2279;
        11'd 934:out = 14'd 2254;
        11'd 935:out = 14'd 2229;
        11'd 936:out = 14'd 2204;
        11'd 937:out = 14'd 2180;
        11'd 938:out = 14'd 2155;
        11'd 939:out = 14'd 2130;
        11'd 940:out = 14'd 2105;
        11'd 941:out = 14'd 2080;
        11'd 942:out = 14'd 2055;
        11'd 943:out = 14'd 2030;
        11'd 944:out = 14'd 2005;
        11'd 945:out = 14'd 1980;
        11'd 946:out = 14'd 1955;
        11'd 947:out = 14'd 1930;
        11'd 948:out = 14'd 1905;
        11'd 949:out = 14'd 1880;
        11'd 950:out = 14'd 1855;
        11'd 951:out = 14'd 1830;
        11'd 952:out = 14'd 1805;
        11'd 953:out = 14'd 1780;
        11'd 954:out = 14'd 1755;
        11'd 955:out = 14'd 1730;
        11'd 956:out = 14'd 1705;
        11'd 957:out = 14'd 1680;
        11'd 958:out = 14'd 1655;
        11'd 959:out = 14'd 1630;
        11'd 960:out = 14'd 1605;
        11'd 961:out = 14'd 1580;
        11'd 962:out = 14'd 1555;
        11'd 963:out = 14'd 1530;
        11'd 964:out = 14'd 1505;
        11'd 965:out = 14'd 1480;
        11'd 966:out = 14'd 1455;
        11'd 967:out = 14'd 1430;
        11'd 968:out = 14'd 1405;
        11'd 969:out = 14'd 1380;
        11'd 970:out = 14'd 1355;
        11'd 971:out = 14'd 1330;
        11'd 972:out = 14'd 1305;
        11'd 973:out = 14'd 1280;
        11'd 974:out = 14'd 1255;
        11'd 975:out = 14'd 1230;
        11'd 976:out = 14'd 1205;
        11'd 977:out = 14'd 1180;
        11'd 978:out = 14'd 1155;
        11'd 979:out = 14'd 1130;
        11'd 980:out = 14'd 1105;
        11'd 981:out = 14'd 1079;
        11'd 982:out = 14'd 1054;
        11'd 983:out = 14'd 1029;
        11'd 984:out = 14'd 1004;
        11'd 985:out = 14'd 979;
        11'd 986:out = 14'd 954;
        11'd 987:out = 14'd 929;
        11'd 988:out = 14'd 904;
        11'd 989:out = 14'd 879;
        11'd 990:out = 14'd 854;
        11'd 991:out = 14'd 829;
        11'd 992:out = 14'd 803;
        11'd 993:out = 14'd 778;
        11'd 994:out = 14'd 753;
        11'd 995:out = 14'd 728;
        11'd 996:out = 14'd 703;
        11'd 997:out = 14'd 678;
        11'd 998:out = 14'd 653;
        11'd 999:out = 14'd 628;
        11'd 1000:out = 14'd 603;
        11'd 1001:out = 14'd 577;
        11'd 1002:out = 14'd 552;
        11'd 1003:out = 14'd 527;
        11'd 1004:out = 14'd 502;
        11'd 1005:out = 14'd 477;
        11'd 1006:out = 14'd 452;
        11'd 1007:out = 14'd 427;
        11'd 1008:out = 14'd 402;
        11'd 1009:out = 14'd 376;
        11'd 1010:out = 14'd 351;
        11'd 1011:out = 14'd 326;
        11'd 1012:out = 14'd 301;
        11'd 1013:out = 14'd 276;
        11'd 1014:out = 14'd 251;
        11'd 1015:out = 14'd 226;
        11'd 1016:out = 14'd 201;
        11'd 1017:out = 14'd 175;
        11'd 1018:out = 14'd 150;
        11'd 1019:out = 14'd 125;
        11'd 1020:out = 14'd 100;
        11'd 1021:out = 14'd 75;
        11'd 1022:out = 14'd 50;
        11'd 1023:out = 14'd 25;
        default: out = 14'd0;
        endcase
    end
    
endmodule
