
module Decoder(
input clk,
input rst,
// 解调结束
input demodulation_down_to_decoder,
// 接收到解调结束信号
output reg demodulation_to_decoder_receive,
// 解调后的数据
input [1535:0] initial_value_input,
// 初始比特流
input [255:0] demodulation_prototype_sequence,
// 输出初始的信息序列
output reg [255:0] prototype_sequence,
// 译码过后的信息序列，用于计算误比特率
output reg [255:0] decision_information,
// 本次译码结束
output reg decoder_down
);
// 对initial_value进行拆分
wire [5:0] initial_value[255:0];
assign initial_value[0] = initial_value_input[5:0];
assign initial_value[1] = initial_value_input[11:6];
assign initial_value[2] = initial_value_input[17:12];
assign initial_value[3] = initial_value_input[23:18];
assign initial_value[4] = initial_value_input[29:24];
assign initial_value[5] = initial_value_input[35:30];
assign initial_value[6] = initial_value_input[41:36];
assign initial_value[7] = initial_value_input[47:42];
assign initial_value[8] = initial_value_input[53:48];
assign initial_value[9] = initial_value_input[59:54];
assign initial_value[10] = initial_value_input[65:60];
assign initial_value[11] = initial_value_input[71:66];
assign initial_value[12] = initial_value_input[77:72];
assign initial_value[13] = initial_value_input[83:78];
assign initial_value[14] = initial_value_input[89:84];
assign initial_value[15] = initial_value_input[95:90];
assign initial_value[16] = initial_value_input[101:96];
assign initial_value[17] = initial_value_input[107:102];
assign initial_value[18] = initial_value_input[113:108];
assign initial_value[19] = initial_value_input[119:114];
assign initial_value[20] = initial_value_input[125:120];
assign initial_value[21] = initial_value_input[131:126];
assign initial_value[22] = initial_value_input[137:132];
assign initial_value[23] = initial_value_input[143:138];
assign initial_value[24] = initial_value_input[149:144];
assign initial_value[25] = initial_value_input[155:150];
assign initial_value[26] = initial_value_input[161:156];
assign initial_value[27] = initial_value_input[167:162];
assign initial_value[28] = initial_value_input[173:168];
assign initial_value[29] = initial_value_input[179:174];
assign initial_value[30] = initial_value_input[185:180];
assign initial_value[31] = initial_value_input[191:186];
assign initial_value[32] = initial_value_input[197:192];
assign initial_value[33] = initial_value_input[203:198];
assign initial_value[34] = initial_value_input[209:204];
assign initial_value[35] = initial_value_input[215:210];
assign initial_value[36] = initial_value_input[221:216];
assign initial_value[37] = initial_value_input[227:222];
assign initial_value[38] = initial_value_input[233:228];
assign initial_value[39] = initial_value_input[239:234];
assign initial_value[40] = initial_value_input[245:240];
assign initial_value[41] = initial_value_input[251:246];
assign initial_value[42] = initial_value_input[257:252];
assign initial_value[43] = initial_value_input[263:258];
assign initial_value[44] = initial_value_input[269:264];
assign initial_value[45] = initial_value_input[275:270];
assign initial_value[46] = initial_value_input[281:276];
assign initial_value[47] = initial_value_input[287:282];
assign initial_value[48] = initial_value_input[293:288];
assign initial_value[49] = initial_value_input[299:294];
assign initial_value[50] = initial_value_input[305:300];
assign initial_value[51] = initial_value_input[311:306];
assign initial_value[52] = initial_value_input[317:312];
assign initial_value[53] = initial_value_input[323:318];
assign initial_value[54] = initial_value_input[329:324];
assign initial_value[55] = initial_value_input[335:330];
assign initial_value[56] = initial_value_input[341:336];
assign initial_value[57] = initial_value_input[347:342];
assign initial_value[58] = initial_value_input[353:348];
assign initial_value[59] = initial_value_input[359:354];
assign initial_value[60] = initial_value_input[365:360];
assign initial_value[61] = initial_value_input[371:366];
assign initial_value[62] = initial_value_input[377:372];
assign initial_value[63] = initial_value_input[383:378];
assign initial_value[64] = initial_value_input[389:384];
assign initial_value[65] = initial_value_input[395:390];
assign initial_value[66] = initial_value_input[401:396];
assign initial_value[67] = initial_value_input[407:402];
assign initial_value[68] = initial_value_input[413:408];
assign initial_value[69] = initial_value_input[419:414];
assign initial_value[70] = initial_value_input[425:420];
assign initial_value[71] = initial_value_input[431:426];
assign initial_value[72] = initial_value_input[437:432];
assign initial_value[73] = initial_value_input[443:438];
assign initial_value[74] = initial_value_input[449:444];
assign initial_value[75] = initial_value_input[455:450];
assign initial_value[76] = initial_value_input[461:456];
assign initial_value[77] = initial_value_input[467:462];
assign initial_value[78] = initial_value_input[473:468];
assign initial_value[79] = initial_value_input[479:474];
assign initial_value[80] = initial_value_input[485:480];
assign initial_value[81] = initial_value_input[491:486];
assign initial_value[82] = initial_value_input[497:492];
assign initial_value[83] = initial_value_input[503:498];
assign initial_value[84] = initial_value_input[509:504];
assign initial_value[85] = initial_value_input[515:510];
assign initial_value[86] = initial_value_input[521:516];
assign initial_value[87] = initial_value_input[527:522];
assign initial_value[88] = initial_value_input[533:528];
assign initial_value[89] = initial_value_input[539:534];
assign initial_value[90] = initial_value_input[545:540];
assign initial_value[91] = initial_value_input[551:546];
assign initial_value[92] = initial_value_input[557:552];
assign initial_value[93] = initial_value_input[563:558];
assign initial_value[94] = initial_value_input[569:564];
assign initial_value[95] = initial_value_input[575:570];
assign initial_value[96] = initial_value_input[581:576];
assign initial_value[97] = initial_value_input[587:582];
assign initial_value[98] = initial_value_input[593:588];
assign initial_value[99] = initial_value_input[599:594];
assign initial_value[100] = initial_value_input[605:600];
assign initial_value[101] = initial_value_input[611:606];
assign initial_value[102] = initial_value_input[617:612];
assign initial_value[103] = initial_value_input[623:618];
assign initial_value[104] = initial_value_input[629:624];
assign initial_value[105] = initial_value_input[635:630];
assign initial_value[106] = initial_value_input[641:636];
assign initial_value[107] = initial_value_input[647:642];
assign initial_value[108] = initial_value_input[653:648];
assign initial_value[109] = initial_value_input[659:654];
assign initial_value[110] = initial_value_input[665:660];
assign initial_value[111] = initial_value_input[671:666];
assign initial_value[112] = initial_value_input[677:672];
assign initial_value[113] = initial_value_input[683:678];
assign initial_value[114] = initial_value_input[689:684];
assign initial_value[115] = initial_value_input[695:690];
assign initial_value[116] = initial_value_input[701:696];
assign initial_value[117] = initial_value_input[707:702];
assign initial_value[118] = initial_value_input[713:708];
assign initial_value[119] = initial_value_input[719:714];
assign initial_value[120] = initial_value_input[725:720];
assign initial_value[121] = initial_value_input[731:726];
assign initial_value[122] = initial_value_input[737:732];
assign initial_value[123] = initial_value_input[743:738];
assign initial_value[124] = initial_value_input[749:744];
assign initial_value[125] = initial_value_input[755:750];
assign initial_value[126] = initial_value_input[761:756];
assign initial_value[127] = initial_value_input[767:762];
assign initial_value[128] = initial_value_input[773:768];
assign initial_value[129] = initial_value_input[779:774];
assign initial_value[130] = initial_value_input[785:780];
assign initial_value[131] = initial_value_input[791:786];
assign initial_value[132] = initial_value_input[797:792];
assign initial_value[133] = initial_value_input[803:798];
assign initial_value[134] = initial_value_input[809:804];
assign initial_value[135] = initial_value_input[815:810];
assign initial_value[136] = initial_value_input[821:816];
assign initial_value[137] = initial_value_input[827:822];
assign initial_value[138] = initial_value_input[833:828];
assign initial_value[139] = initial_value_input[839:834];
assign initial_value[140] = initial_value_input[845:840];
assign initial_value[141] = initial_value_input[851:846];
assign initial_value[142] = initial_value_input[857:852];
assign initial_value[143] = initial_value_input[863:858];
assign initial_value[144] = initial_value_input[869:864];
assign initial_value[145] = initial_value_input[875:870];
assign initial_value[146] = initial_value_input[881:876];
assign initial_value[147] = initial_value_input[887:882];
assign initial_value[148] = initial_value_input[893:888];
assign initial_value[149] = initial_value_input[899:894];
assign initial_value[150] = initial_value_input[905:900];
assign initial_value[151] = initial_value_input[911:906];
assign initial_value[152] = initial_value_input[917:912];
assign initial_value[153] = initial_value_input[923:918];
assign initial_value[154] = initial_value_input[929:924];
assign initial_value[155] = initial_value_input[935:930];
assign initial_value[156] = initial_value_input[941:936];
assign initial_value[157] = initial_value_input[947:942];
assign initial_value[158] = initial_value_input[953:948];
assign initial_value[159] = initial_value_input[959:954];
assign initial_value[160] = initial_value_input[965:960];
assign initial_value[161] = initial_value_input[971:966];
assign initial_value[162] = initial_value_input[977:972];
assign initial_value[163] = initial_value_input[983:978];
assign initial_value[164] = initial_value_input[989:984];
assign initial_value[165] = initial_value_input[995:990];
assign initial_value[166] = initial_value_input[1001:996];
assign initial_value[167] = initial_value_input[1007:1002];
assign initial_value[168] = initial_value_input[1013:1008];
assign initial_value[169] = initial_value_input[1019:1014];
assign initial_value[170] = initial_value_input[1025:1020];
assign initial_value[171] = initial_value_input[1031:1026];
assign initial_value[172] = initial_value_input[1037:1032];
assign initial_value[173] = initial_value_input[1043:1038];
assign initial_value[174] = initial_value_input[1049:1044];
assign initial_value[175] = initial_value_input[1055:1050];
assign initial_value[176] = initial_value_input[1061:1056];
assign initial_value[177] = initial_value_input[1067:1062];
assign initial_value[178] = initial_value_input[1073:1068];
assign initial_value[179] = initial_value_input[1079:1074];
assign initial_value[180] = initial_value_input[1085:1080];
assign initial_value[181] = initial_value_input[1091:1086];
assign initial_value[182] = initial_value_input[1097:1092];
assign initial_value[183] = initial_value_input[1103:1098];
assign initial_value[184] = initial_value_input[1109:1104];
assign initial_value[185] = initial_value_input[1115:1110];
assign initial_value[186] = initial_value_input[1121:1116];
assign initial_value[187] = initial_value_input[1127:1122];
assign initial_value[188] = initial_value_input[1133:1128];
assign initial_value[189] = initial_value_input[1139:1134];
assign initial_value[190] = initial_value_input[1145:1140];
assign initial_value[191] = initial_value_input[1151:1146];
assign initial_value[192] = initial_value_input[1157:1152];
assign initial_value[193] = initial_value_input[1163:1158];
assign initial_value[194] = initial_value_input[1169:1164];
assign initial_value[195] = initial_value_input[1175:1170];
assign initial_value[196] = initial_value_input[1181:1176];
assign initial_value[197] = initial_value_input[1187:1182];
assign initial_value[198] = initial_value_input[1193:1188];
assign initial_value[199] = initial_value_input[1199:1194];
assign initial_value[200] = initial_value_input[1205:1200];
assign initial_value[201] = initial_value_input[1211:1206];
assign initial_value[202] = initial_value_input[1217:1212];
assign initial_value[203] = initial_value_input[1223:1218];
assign initial_value[204] = initial_value_input[1229:1224];
assign initial_value[205] = initial_value_input[1235:1230];
assign initial_value[206] = initial_value_input[1241:1236];
assign initial_value[207] = initial_value_input[1247:1242];
assign initial_value[208] = initial_value_input[1253:1248];
assign initial_value[209] = initial_value_input[1259:1254];
assign initial_value[210] = initial_value_input[1265:1260];
assign initial_value[211] = initial_value_input[1271:1266];
assign initial_value[212] = initial_value_input[1277:1272];
assign initial_value[213] = initial_value_input[1283:1278];
assign initial_value[214] = initial_value_input[1289:1284];
assign initial_value[215] = initial_value_input[1295:1290];
assign initial_value[216] = initial_value_input[1301:1296];
assign initial_value[217] = initial_value_input[1307:1302];
assign initial_value[218] = initial_value_input[1313:1308];
assign initial_value[219] = initial_value_input[1319:1314];
assign initial_value[220] = initial_value_input[1325:1320];
assign initial_value[221] = initial_value_input[1331:1326];
assign initial_value[222] = initial_value_input[1337:1332];
assign initial_value[223] = initial_value_input[1343:1338];
assign initial_value[224] = initial_value_input[1349:1344];
assign initial_value[225] = initial_value_input[1355:1350];
assign initial_value[226] = initial_value_input[1361:1356];
assign initial_value[227] = initial_value_input[1367:1362];
assign initial_value[228] = initial_value_input[1373:1368];
assign initial_value[229] = initial_value_input[1379:1374];
assign initial_value[230] = initial_value_input[1385:1380];
assign initial_value[231] = initial_value_input[1391:1386];
assign initial_value[232] = initial_value_input[1397:1392];
assign initial_value[233] = initial_value_input[1403:1398];
assign initial_value[234] = initial_value_input[1409:1404];
assign initial_value[235] = initial_value_input[1415:1410];
assign initial_value[236] = initial_value_input[1421:1416];
assign initial_value[237] = initial_value_input[1427:1422];
assign initial_value[238] = initial_value_input[1433:1428];
assign initial_value[239] = initial_value_input[1439:1434];
assign initial_value[240] = initial_value_input[1445:1440];
assign initial_value[241] = initial_value_input[1451:1446];
assign initial_value[242] = initial_value_input[1457:1452];
assign initial_value[243] = initial_value_input[1463:1458];
assign initial_value[244] = initial_value_input[1469:1464];
assign initial_value[245] = initial_value_input[1475:1470];
assign initial_value[246] = initial_value_input[1481:1476];
assign initial_value[247] = initial_value_input[1487:1482];
assign initial_value[248] = initial_value_input[1493:1488];
assign initial_value[249] = initial_value_input[1499:1494];
assign initial_value[250] = initial_value_input[1505:1500];
assign initial_value[251] = initial_value_input[1511:1506];
assign initial_value[252] = initial_value_input[1517:1512];
assign initial_value[253] = initial_value_input[1523:1518];
assign initial_value[254] = initial_value_input[1529:1524];
assign initial_value[255] = initial_value_input[1535:1530];


// 定义跟判决部分有关的变量
reg [255:0]initial_value_enable;
wire [255:0]initial_down;
reg check_begin;
reg [2:0] decision_state;
reg decision_down;
reg decision_success;
reg [9:0] decision_times;
reg [255:0]decision_result;
reg decision_time_max;
wire [255:0]decision_variable_enable;


// 校验节点0的接口
wire [35:0] value_variable_to_check_0;
wire [35:0] value_check_0_to_variable;
wire [5:0] enable_variable_to_check_0;
wire [5:0] enable_check_0_to_variable;

// 拆分后校验节点0传递给变量节点0的值以及对变量节点0传递过来的值
wire [5:0] value_check_0_to_variable_0;
wire enable_check_0_to_variable_0;
wire [5:0] value_variable_0_to_check_0;
wire enable_variable_0_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_0 = value_check_0_to_variable[5:0];
assign enable_check_0_to_variable_0 = enable_check_0_to_variable[0];
// 对变量节点0传递过来的值进行组合
assign value_variable_to_check_0[5:0] = value_variable_0_to_check_0;
assign enable_variable_to_check_0[0] = enable_variable_0_to_check_0;

// 拆分后校验节点0传递给变量节点43的值以及对变量节点43传递过来的值
wire [5:0] value_check_0_to_variable_43;
wire enable_check_0_to_variable_43;
wire [5:0] value_variable_43_to_check_0;
wire enable_variable_43_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_43 = value_check_0_to_variable[11:6];
assign enable_check_0_to_variable_43 = enable_check_0_to_variable[1];
// 对变量节点43传递过来的值进行组合
assign value_variable_to_check_0[11:6] = value_variable_43_to_check_0;
assign enable_variable_to_check_0[1] = enable_variable_43_to_check_0;

// 拆分后校验节点0传递给变量节点86的值以及对变量节点86传递过来的值
wire [5:0] value_check_0_to_variable_86;
wire enable_check_0_to_variable_86;
wire [5:0] value_variable_86_to_check_0;
wire enable_variable_86_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_86 = value_check_0_to_variable[17:12];
assign enable_check_0_to_variable_86 = enable_check_0_to_variable[2];
// 对变量节点86传递过来的值进行组合
assign value_variable_to_check_0[17:12] = value_variable_86_to_check_0;
assign enable_variable_to_check_0[2] = enable_variable_86_to_check_0;

// 拆分后校验节点0传递给变量节点131的值以及对变量节点131传递过来的值
wire [5:0] value_check_0_to_variable_131;
wire enable_check_0_to_variable_131;
wire [5:0] value_variable_131_to_check_0;
wire enable_variable_131_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_131 = value_check_0_to_variable[23:18];
assign enable_check_0_to_variable_131 = enable_check_0_to_variable[3];
// 对变量节点131传递过来的值进行组合
assign value_variable_to_check_0[23:18] = value_variable_131_to_check_0;
assign enable_variable_to_check_0[3] = enable_variable_131_to_check_0;

// 拆分后校验节点0传递给变量节点170的值以及对变量节点170传递过来的值
wire [5:0] value_check_0_to_variable_170;
wire enable_check_0_to_variable_170;
wire [5:0] value_variable_170_to_check_0;
wire enable_variable_170_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_170 = value_check_0_to_variable[29:24];
assign enable_check_0_to_variable_170 = enable_check_0_to_variable[4];
// 对变量节点170传递过来的值进行组合
assign value_variable_to_check_0[29:24] = value_variable_170_to_check_0;
assign enable_variable_to_check_0[4] = enable_variable_170_to_check_0;

// 拆分后校验节点0传递给变量节点214的值以及对变量节点214传递过来的值
wire [5:0] value_check_0_to_variable_214;
wire enable_check_0_to_variable_214;
wire [5:0] value_variable_214_to_check_0;
wire enable_variable_214_to_check_0;
// 对校验节点0的输出值进行拆分
assign value_check_0_to_variable_214 = value_check_0_to_variable[35:30];
assign enable_check_0_to_variable_214 = enable_check_0_to_variable[5];
// 对变量节点214传递过来的值进行组合
assign value_variable_to_check_0[35:30] = value_variable_214_to_check_0;
assign enable_variable_to_check_0[5] = enable_variable_214_to_check_0;


// 校验节点1的接口
wire [35:0] value_variable_to_check_1;
wire [35:0] value_check_1_to_variable;
wire [5:0] enable_variable_to_check_1;
wire [5:0] enable_check_1_to_variable;

// 拆分后校验节点1传递给变量节点1的值以及对变量节点1传递过来的值
wire [5:0] value_check_1_to_variable_1;
wire enable_check_1_to_variable_1;
wire [5:0] value_variable_1_to_check_1;
wire enable_variable_1_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_1 = value_check_1_to_variable[5:0];
assign enable_check_1_to_variable_1 = enable_check_1_to_variable[0];
// 对变量节点1传递过来的值进行组合
assign value_variable_to_check_1[5:0] = value_variable_1_to_check_1;
assign enable_variable_to_check_1[0] = enable_variable_1_to_check_1;

// 拆分后校验节点1传递给变量节点42的值以及对变量节点42传递过来的值
wire [5:0] value_check_1_to_variable_42;
wire enable_check_1_to_variable_42;
wire [5:0] value_variable_42_to_check_1;
wire enable_variable_42_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_42 = value_check_1_to_variable[11:6];
assign enable_check_1_to_variable_42 = enable_check_1_to_variable[1];
// 对变量节点42传递过来的值进行组合
assign value_variable_to_check_1[11:6] = value_variable_42_to_check_1;
assign enable_variable_to_check_1[1] = enable_variable_42_to_check_1;

// 拆分后校验节点1传递给变量节点87的值以及对变量节点87传递过来的值
wire [5:0] value_check_1_to_variable_87;
wire enable_check_1_to_variable_87;
wire [5:0] value_variable_87_to_check_1;
wire enable_variable_87_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_87 = value_check_1_to_variable[17:12];
assign enable_check_1_to_variable_87 = enable_check_1_to_variable[2];
// 对变量节点87传递过来的值进行组合
assign value_variable_to_check_1[17:12] = value_variable_87_to_check_1;
assign enable_variable_to_check_1[2] = enable_variable_87_to_check_1;

// 拆分后校验节点1传递给变量节点132的值以及对变量节点132传递过来的值
wire [5:0] value_check_1_to_variable_132;
wire enable_check_1_to_variable_132;
wire [5:0] value_variable_132_to_check_1;
wire enable_variable_132_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_132 = value_check_1_to_variable[23:18];
assign enable_check_1_to_variable_132 = enable_check_1_to_variable[3];
// 对变量节点132传递过来的值进行组合
assign value_variable_to_check_1[23:18] = value_variable_132_to_check_1;
assign enable_variable_to_check_1[3] = enable_variable_132_to_check_1;

// 拆分后校验节点1传递给变量节点173的值以及对变量节点173传递过来的值
wire [5:0] value_check_1_to_variable_173;
wire enable_check_1_to_variable_173;
wire [5:0] value_variable_173_to_check_1;
wire enable_variable_173_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_173 = value_check_1_to_variable[29:24];
assign enable_check_1_to_variable_173 = enable_check_1_to_variable[4];
// 对变量节点173传递过来的值进行组合
assign value_variable_to_check_1[29:24] = value_variable_173_to_check_1;
assign enable_variable_to_check_1[4] = enable_variable_173_to_check_1;

// 拆分后校验节点1传递给变量节点215的值以及对变量节点215传递过来的值
wire [5:0] value_check_1_to_variable_215;
wire enable_check_1_to_variable_215;
wire [5:0] value_variable_215_to_check_1;
wire enable_variable_215_to_check_1;
// 对校验节点1的输出值进行拆分
assign value_check_1_to_variable_215 = value_check_1_to_variable[35:30];
assign enable_check_1_to_variable_215 = enable_check_1_to_variable[5];
// 对变量节点215传递过来的值进行组合
assign value_variable_to_check_1[35:30] = value_variable_215_to_check_1;
assign enable_variable_to_check_1[5] = enable_variable_215_to_check_1;


// 校验节点2的接口
wire [35:0] value_variable_to_check_2;
wire [35:0] value_check_2_to_variable;
wire [5:0] enable_variable_to_check_2;
wire [5:0] enable_check_2_to_variable;

// 拆分后校验节点2传递给变量节点2的值以及对变量节点2传递过来的值
wire [5:0] value_check_2_to_variable_2;
wire enable_check_2_to_variable_2;
wire [5:0] value_variable_2_to_check_2;
wire enable_variable_2_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_2 = value_check_2_to_variable[5:0];
assign enable_check_2_to_variable_2 = enable_check_2_to_variable[0];
// 对变量节点2传递过来的值进行组合
assign value_variable_to_check_2[5:0] = value_variable_2_to_check_2;
assign enable_variable_to_check_2[0] = enable_variable_2_to_check_2;

// 拆分后校验节点2传递给变量节点44的值以及对变量节点44传递过来的值
wire [5:0] value_check_2_to_variable_44;
wire enable_check_2_to_variable_44;
wire [5:0] value_variable_44_to_check_2;
wire enable_variable_44_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_44 = value_check_2_to_variable[11:6];
assign enable_check_2_to_variable_44 = enable_check_2_to_variable[1];
// 对变量节点44传递过来的值进行组合
assign value_variable_to_check_2[11:6] = value_variable_44_to_check_2;
assign enable_variable_to_check_2[1] = enable_variable_44_to_check_2;

// 拆分后校验节点2传递给变量节点88的值以及对变量节点88传递过来的值
wire [5:0] value_check_2_to_variable_88;
wire enable_check_2_to_variable_88;
wire [5:0] value_variable_88_to_check_2;
wire enable_variable_88_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_88 = value_check_2_to_variable[17:12];
assign enable_check_2_to_variable_88 = enable_check_2_to_variable[2];
// 对变量节点88传递过来的值进行组合
assign value_variable_to_check_2[17:12] = value_variable_88_to_check_2;
assign enable_variable_to_check_2[2] = enable_variable_88_to_check_2;

// 拆分后校验节点2传递给变量节点133的值以及对变量节点133传递过来的值
wire [5:0] value_check_2_to_variable_133;
wire enable_check_2_to_variable_133;
wire [5:0] value_variable_133_to_check_2;
wire enable_variable_133_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_133 = value_check_2_to_variable[23:18];
assign enable_check_2_to_variable_133 = enable_check_2_to_variable[3];
// 对变量节点133传递过来的值进行组合
assign value_variable_to_check_2[23:18] = value_variable_133_to_check_2;
assign enable_variable_to_check_2[3] = enable_variable_133_to_check_2;

// 拆分后校验节点2传递给变量节点174的值以及对变量节点174传递过来的值
wire [5:0] value_check_2_to_variable_174;
wire enable_check_2_to_variable_174;
wire [5:0] value_variable_174_to_check_2;
wire enable_variable_174_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_174 = value_check_2_to_variable[29:24];
assign enable_check_2_to_variable_174 = enable_check_2_to_variable[4];
// 对变量节点174传递过来的值进行组合
assign value_variable_to_check_2[29:24] = value_variable_174_to_check_2;
assign enable_variable_to_check_2[4] = enable_variable_174_to_check_2;

// 拆分后校验节点2传递给变量节点216的值以及对变量节点216传递过来的值
wire [5:0] value_check_2_to_variable_216;
wire enable_check_2_to_variable_216;
wire [5:0] value_variable_216_to_check_2;
wire enable_variable_216_to_check_2;
// 对校验节点2的输出值进行拆分
assign value_check_2_to_variable_216 = value_check_2_to_variable[35:30];
assign enable_check_2_to_variable_216 = enable_check_2_to_variable[5];
// 对变量节点216传递过来的值进行组合
assign value_variable_to_check_2[35:30] = value_variable_216_to_check_2;
assign enable_variable_to_check_2[5] = enable_variable_216_to_check_2;


// 校验节点3的接口
wire [35:0] value_variable_to_check_3;
wire [35:0] value_check_3_to_variable;
wire [5:0] enable_variable_to_check_3;
wire [5:0] enable_check_3_to_variable;

// 拆分后校验节点3传递给变量节点3的值以及对变量节点3传递过来的值
wire [5:0] value_check_3_to_variable_3;
wire enable_check_3_to_variable_3;
wire [5:0] value_variable_3_to_check_3;
wire enable_variable_3_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_3 = value_check_3_to_variable[5:0];
assign enable_check_3_to_variable_3 = enable_check_3_to_variable[0];
// 对变量节点3传递过来的值进行组合
assign value_variable_to_check_3[5:0] = value_variable_3_to_check_3;
assign enable_variable_to_check_3[0] = enable_variable_3_to_check_3;

// 拆分后校验节点3传递给变量节点45的值以及对变量节点45传递过来的值
wire [5:0] value_check_3_to_variable_45;
wire enable_check_3_to_variable_45;
wire [5:0] value_variable_45_to_check_3;
wire enable_variable_45_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_45 = value_check_3_to_variable[11:6];
assign enable_check_3_to_variable_45 = enable_check_3_to_variable[1];
// 对变量节点45传递过来的值进行组合
assign value_variable_to_check_3[11:6] = value_variable_45_to_check_3;
assign enable_variable_to_check_3[1] = enable_variable_45_to_check_3;

// 拆分后校验节点3传递给变量节点89的值以及对变量节点89传递过来的值
wire [5:0] value_check_3_to_variable_89;
wire enable_check_3_to_variable_89;
wire [5:0] value_variable_89_to_check_3;
wire enable_variable_89_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_89 = value_check_3_to_variable[17:12];
assign enable_check_3_to_variable_89 = enable_check_3_to_variable[2];
// 对变量节点89传递过来的值进行组合
assign value_variable_to_check_3[17:12] = value_variable_89_to_check_3;
assign enable_variable_to_check_3[2] = enable_variable_89_to_check_3;

// 拆分后校验节点3传递给变量节点134的值以及对变量节点134传递过来的值
wire [5:0] value_check_3_to_variable_134;
wire enable_check_3_to_variable_134;
wire [5:0] value_variable_134_to_check_3;
wire enable_variable_134_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_134 = value_check_3_to_variable[23:18];
assign enable_check_3_to_variable_134 = enable_check_3_to_variable[3];
// 对变量节点134传递过来的值进行组合
assign value_variable_to_check_3[23:18] = value_variable_134_to_check_3;
assign enable_variable_to_check_3[3] = enable_variable_134_to_check_3;

// 拆分后校验节点3传递给变量节点175的值以及对变量节点175传递过来的值
wire [5:0] value_check_3_to_variable_175;
wire enable_check_3_to_variable_175;
wire [5:0] value_variable_175_to_check_3;
wire enable_variable_175_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_175 = value_check_3_to_variable[29:24];
assign enable_check_3_to_variable_175 = enable_check_3_to_variable[4];
// 对变量节点175传递过来的值进行组合
assign value_variable_to_check_3[29:24] = value_variable_175_to_check_3;
assign enable_variable_to_check_3[4] = enable_variable_175_to_check_3;

// 拆分后校验节点3传递给变量节点217的值以及对变量节点217传递过来的值
wire [5:0] value_check_3_to_variable_217;
wire enable_check_3_to_variable_217;
wire [5:0] value_variable_217_to_check_3;
wire enable_variable_217_to_check_3;
// 对校验节点3的输出值进行拆分
assign value_check_3_to_variable_217 = value_check_3_to_variable[35:30];
assign enable_check_3_to_variable_217 = enable_check_3_to_variable[5];
// 对变量节点217传递过来的值进行组合
assign value_variable_to_check_3[35:30] = value_variable_217_to_check_3;
assign enable_variable_to_check_3[5] = enable_variable_217_to_check_3;


// 校验节点4的接口
wire [35:0] value_variable_to_check_4;
wire [35:0] value_check_4_to_variable;
wire [5:0] enable_variable_to_check_4;
wire [5:0] enable_check_4_to_variable;

// 拆分后校验节点4传递给变量节点4的值以及对变量节点4传递过来的值
wire [5:0] value_check_4_to_variable_4;
wire enable_check_4_to_variable_4;
wire [5:0] value_variable_4_to_check_4;
wire enable_variable_4_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_4 = value_check_4_to_variable[5:0];
assign enable_check_4_to_variable_4 = enable_check_4_to_variable[0];
// 对变量节点4传递过来的值进行组合
assign value_variable_to_check_4[5:0] = value_variable_4_to_check_4;
assign enable_variable_to_check_4[0] = enable_variable_4_to_check_4;

// 拆分后校验节点4传递给变量节点46的值以及对变量节点46传递过来的值
wire [5:0] value_check_4_to_variable_46;
wire enable_check_4_to_variable_46;
wire [5:0] value_variable_46_to_check_4;
wire enable_variable_46_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_46 = value_check_4_to_variable[11:6];
assign enable_check_4_to_variable_46 = enable_check_4_to_variable[1];
// 对变量节点46传递过来的值进行组合
assign value_variable_to_check_4[11:6] = value_variable_46_to_check_4;
assign enable_variable_to_check_4[1] = enable_variable_46_to_check_4;

// 拆分后校验节点4传递给变量节点90的值以及对变量节点90传递过来的值
wire [5:0] value_check_4_to_variable_90;
wire enable_check_4_to_variable_90;
wire [5:0] value_variable_90_to_check_4;
wire enable_variable_90_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_90 = value_check_4_to_variable[17:12];
assign enable_check_4_to_variable_90 = enable_check_4_to_variable[2];
// 对变量节点90传递过来的值进行组合
assign value_variable_to_check_4[17:12] = value_variable_90_to_check_4;
assign enable_variable_to_check_4[2] = enable_variable_90_to_check_4;

// 拆分后校验节点4传递给变量节点128的值以及对变量节点128传递过来的值
wire [5:0] value_check_4_to_variable_128;
wire enable_check_4_to_variable_128;
wire [5:0] value_variable_128_to_check_4;
wire enable_variable_128_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_128 = value_check_4_to_variable[23:18];
assign enable_check_4_to_variable_128 = enable_check_4_to_variable[3];
// 对变量节点128传递过来的值进行组合
assign value_variable_to_check_4[23:18] = value_variable_128_to_check_4;
assign enable_variable_to_check_4[3] = enable_variable_128_to_check_4;

// 拆分后校验节点4传递给变量节点176的值以及对变量节点176传递过来的值
wire [5:0] value_check_4_to_variable_176;
wire enable_check_4_to_variable_176;
wire [5:0] value_variable_176_to_check_4;
wire enable_variable_176_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_176 = value_check_4_to_variable[29:24];
assign enable_check_4_to_variable_176 = enable_check_4_to_variable[4];
// 对变量节点176传递过来的值进行组合
assign value_variable_to_check_4[29:24] = value_variable_176_to_check_4;
assign enable_variable_to_check_4[4] = enable_variable_176_to_check_4;

// 拆分后校验节点4传递给变量节点218的值以及对变量节点218传递过来的值
wire [5:0] value_check_4_to_variable_218;
wire enable_check_4_to_variable_218;
wire [5:0] value_variable_218_to_check_4;
wire enable_variable_218_to_check_4;
// 对校验节点4的输出值进行拆分
assign value_check_4_to_variable_218 = value_check_4_to_variable[35:30];
assign enable_check_4_to_variable_218 = enable_check_4_to_variable[5];
// 对变量节点218传递过来的值进行组合
assign value_variable_to_check_4[35:30] = value_variable_218_to_check_4;
assign enable_variable_to_check_4[5] = enable_variable_218_to_check_4;


// 校验节点5的接口
wire [35:0] value_variable_to_check_5;
wire [35:0] value_check_5_to_variable;
wire [5:0] enable_variable_to_check_5;
wire [5:0] enable_check_5_to_variable;

// 拆分后校验节点5传递给变量节点5的值以及对变量节点5传递过来的值
wire [5:0] value_check_5_to_variable_5;
wire enable_check_5_to_variable_5;
wire [5:0] value_variable_5_to_check_5;
wire enable_variable_5_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_5 = value_check_5_to_variable[5:0];
assign enable_check_5_to_variable_5 = enable_check_5_to_variable[0];
// 对变量节点5传递过来的值进行组合
assign value_variable_to_check_5[5:0] = value_variable_5_to_check_5;
assign enable_variable_to_check_5[0] = enable_variable_5_to_check_5;

// 拆分后校验节点5传递给变量节点47的值以及对变量节点47传递过来的值
wire [5:0] value_check_5_to_variable_47;
wire enable_check_5_to_variable_47;
wire [5:0] value_variable_47_to_check_5;
wire enable_variable_47_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_47 = value_check_5_to_variable[11:6];
assign enable_check_5_to_variable_47 = enable_check_5_to_variable[1];
// 对变量节点47传递过来的值进行组合
assign value_variable_to_check_5[11:6] = value_variable_47_to_check_5;
assign enable_variable_to_check_5[1] = enable_variable_47_to_check_5;

// 拆分后校验节点5传递给变量节点91的值以及对变量节点91传递过来的值
wire [5:0] value_check_5_to_variable_91;
wire enable_check_5_to_variable_91;
wire [5:0] value_variable_91_to_check_5;
wire enable_variable_91_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_91 = value_check_5_to_variable[17:12];
assign enable_check_5_to_variable_91 = enable_check_5_to_variable[2];
// 对变量节点91传递过来的值进行组合
assign value_variable_to_check_5[17:12] = value_variable_91_to_check_5;
assign enable_variable_to_check_5[2] = enable_variable_91_to_check_5;

// 拆分后校验节点5传递给变量节点135的值以及对变量节点135传递过来的值
wire [5:0] value_check_5_to_variable_135;
wire enable_check_5_to_variable_135;
wire [5:0] value_variable_135_to_check_5;
wire enable_variable_135_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_135 = value_check_5_to_variable[23:18];
assign enable_check_5_to_variable_135 = enable_check_5_to_variable[3];
// 对变量节点135传递过来的值进行组合
assign value_variable_to_check_5[23:18] = value_variable_135_to_check_5;
assign enable_variable_to_check_5[3] = enable_variable_135_to_check_5;

// 拆分后校验节点5传递给变量节点177的值以及对变量节点177传递过来的值
wire [5:0] value_check_5_to_variable_177;
wire enable_check_5_to_variable_177;
wire [5:0] value_variable_177_to_check_5;
wire enable_variable_177_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_177 = value_check_5_to_variable[29:24];
assign enable_check_5_to_variable_177 = enable_check_5_to_variable[4];
// 对变量节点177传递过来的值进行组合
assign value_variable_to_check_5[29:24] = value_variable_177_to_check_5;
assign enable_variable_to_check_5[4] = enable_variable_177_to_check_5;

// 拆分后校验节点5传递给变量节点219的值以及对变量节点219传递过来的值
wire [5:0] value_check_5_to_variable_219;
wire enable_check_5_to_variable_219;
wire [5:0] value_variable_219_to_check_5;
wire enable_variable_219_to_check_5;
// 对校验节点5的输出值进行拆分
assign value_check_5_to_variable_219 = value_check_5_to_variable[35:30];
assign enable_check_5_to_variable_219 = enable_check_5_to_variable[5];
// 对变量节点219传递过来的值进行组合
assign value_variable_to_check_5[35:30] = value_variable_219_to_check_5;
assign enable_variable_to_check_5[5] = enable_variable_219_to_check_5;


// 校验节点6的接口
wire [35:0] value_variable_to_check_6;
wire [35:0] value_check_6_to_variable;
wire [5:0] enable_variable_to_check_6;
wire [5:0] enable_check_6_to_variable;

// 拆分后校验节点6传递给变量节点1的值以及对变量节点1传递过来的值
wire [5:0] value_check_6_to_variable_1;
wire enable_check_6_to_variable_1;
wire [5:0] value_variable_1_to_check_6;
wire enable_variable_1_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_1 = value_check_6_to_variable[5:0];
assign enable_check_6_to_variable_1 = enable_check_6_to_variable[0];
// 对变量节点1传递过来的值进行组合
assign value_variable_to_check_6[5:0] = value_variable_1_to_check_6;
assign enable_variable_to_check_6[0] = enable_variable_1_to_check_6;

// 拆分后校验节点6传递给变量节点48的值以及对变量节点48传递过来的值
wire [5:0] value_check_6_to_variable_48;
wire enable_check_6_to_variable_48;
wire [5:0] value_variable_48_to_check_6;
wire enable_variable_48_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_48 = value_check_6_to_variable[11:6];
assign enable_check_6_to_variable_48 = enable_check_6_to_variable[1];
// 对变量节点48传递过来的值进行组合
assign value_variable_to_check_6[11:6] = value_variable_48_to_check_6;
assign enable_variable_to_check_6[1] = enable_variable_48_to_check_6;

// 拆分后校验节点6传递给变量节点92的值以及对变量节点92传递过来的值
wire [5:0] value_check_6_to_variable_92;
wire enable_check_6_to_variable_92;
wire [5:0] value_variable_92_to_check_6;
wire enable_variable_92_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_92 = value_check_6_to_variable[17:12];
assign enable_check_6_to_variable_92 = enable_check_6_to_variable[2];
// 对变量节点92传递过来的值进行组合
assign value_variable_to_check_6[17:12] = value_variable_92_to_check_6;
assign enable_variable_to_check_6[2] = enable_variable_92_to_check_6;

// 拆分后校验节点6传递给变量节点131的值以及对变量节点131传递过来的值
wire [5:0] value_check_6_to_variable_131;
wire enable_check_6_to_variable_131;
wire [5:0] value_variable_131_to_check_6;
wire enable_variable_131_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_131 = value_check_6_to_variable[23:18];
assign enable_check_6_to_variable_131 = enable_check_6_to_variable[3];
// 对变量节点131传递过来的值进行组合
assign value_variable_to_check_6[23:18] = value_variable_131_to_check_6;
assign enable_variable_to_check_6[3] = enable_variable_131_to_check_6;

// 拆分后校验节点6传递给变量节点178的值以及对变量节点178传递过来的值
wire [5:0] value_check_6_to_variable_178;
wire enable_check_6_to_variable_178;
wire [5:0] value_variable_178_to_check_6;
wire enable_variable_178_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_178 = value_check_6_to_variable[29:24];
assign enable_check_6_to_variable_178 = enable_check_6_to_variable[4];
// 对变量节点178传递过来的值进行组合
assign value_variable_to_check_6[29:24] = value_variable_178_to_check_6;
assign enable_variable_to_check_6[4] = enable_variable_178_to_check_6;

// 拆分后校验节点6传递给变量节点220的值以及对变量节点220传递过来的值
wire [5:0] value_check_6_to_variable_220;
wire enable_check_6_to_variable_220;
wire [5:0] value_variable_220_to_check_6;
wire enable_variable_220_to_check_6;
// 对校验节点6的输出值进行拆分
assign value_check_6_to_variable_220 = value_check_6_to_variable[35:30];
assign enable_check_6_to_variable_220 = enable_check_6_to_variable[5];
// 对变量节点220传递过来的值进行组合
assign value_variable_to_check_6[35:30] = value_variable_220_to_check_6;
assign enable_variable_to_check_6[5] = enable_variable_220_to_check_6;


// 校验节点7的接口
wire [35:0] value_variable_to_check_7;
wire [35:0] value_check_7_to_variable;
wire [5:0] enable_variable_to_check_7;
wire [5:0] enable_check_7_to_variable;

// 拆分后校验节点7传递给变量节点6的值以及对变量节点6传递过来的值
wire [5:0] value_check_7_to_variable_6;
wire enable_check_7_to_variable_6;
wire [5:0] value_variable_6_to_check_7;
wire enable_variable_6_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_6 = value_check_7_to_variable[5:0];
assign enable_check_7_to_variable_6 = enable_check_7_to_variable[0];
// 对变量节点6传递过来的值进行组合
assign value_variable_to_check_7[5:0] = value_variable_6_to_check_7;
assign enable_variable_to_check_7[0] = enable_variable_6_to_check_7;

// 拆分后校验节点7传递给变量节点47的值以及对变量节点47传递过来的值
wire [5:0] value_check_7_to_variable_47;
wire enable_check_7_to_variable_47;
wire [5:0] value_variable_47_to_check_7;
wire enable_variable_47_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_47 = value_check_7_to_variable[11:6];
assign enable_check_7_to_variable_47 = enable_check_7_to_variable[1];
// 对变量节点47传递过来的值进行组合
assign value_variable_to_check_7[11:6] = value_variable_47_to_check_7;
assign enable_variable_to_check_7[1] = enable_variable_47_to_check_7;

// 拆分后校验节点7传递给变量节点93的值以及对变量节点93传递过来的值
wire [5:0] value_check_7_to_variable_93;
wire enable_check_7_to_variable_93;
wire [5:0] value_variable_93_to_check_7;
wire enable_variable_93_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_93 = value_check_7_to_variable[17:12];
assign enable_check_7_to_variable_93 = enable_check_7_to_variable[2];
// 对变量节点93传递过来的值进行组合
assign value_variable_to_check_7[17:12] = value_variable_93_to_check_7;
assign enable_variable_to_check_7[2] = enable_variable_93_to_check_7;

// 拆分后校验节点7传递给变量节点136的值以及对变量节点136传递过来的值
wire [5:0] value_check_7_to_variable_136;
wire enable_check_7_to_variable_136;
wire [5:0] value_variable_136_to_check_7;
wire enable_variable_136_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_136 = value_check_7_to_variable[23:18];
assign enable_check_7_to_variable_136 = enable_check_7_to_variable[3];
// 对变量节点136传递过来的值进行组合
assign value_variable_to_check_7[23:18] = value_variable_136_to_check_7;
assign enable_variable_to_check_7[3] = enable_variable_136_to_check_7;

// 拆分后校验节点7传递给变量节点179的值以及对变量节点179传递过来的值
wire [5:0] value_check_7_to_variable_179;
wire enable_check_7_to_variable_179;
wire [5:0] value_variable_179_to_check_7;
wire enable_variable_179_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_179 = value_check_7_to_variable[29:24];
assign enable_check_7_to_variable_179 = enable_check_7_to_variable[4];
// 对变量节点179传递过来的值进行组合
assign value_variable_to_check_7[29:24] = value_variable_179_to_check_7;
assign enable_variable_to_check_7[4] = enable_variable_179_to_check_7;

// 拆分后校验节点7传递给变量节点221的值以及对变量节点221传递过来的值
wire [5:0] value_check_7_to_variable_221;
wire enable_check_7_to_variable_221;
wire [5:0] value_variable_221_to_check_7;
wire enable_variable_221_to_check_7;
// 对校验节点7的输出值进行拆分
assign value_check_7_to_variable_221 = value_check_7_to_variable[35:30];
assign enable_check_7_to_variable_221 = enable_check_7_to_variable[5];
// 对变量节点221传递过来的值进行组合
assign value_variable_to_check_7[35:30] = value_variable_221_to_check_7;
assign enable_variable_to_check_7[5] = enable_variable_221_to_check_7;


// 校验节点8的接口
wire [35:0] value_variable_to_check_8;
wire [35:0] value_check_8_to_variable;
wire [5:0] enable_variable_to_check_8;
wire [5:0] enable_check_8_to_variable;

// 拆分后校验节点8传递给变量节点7的值以及对变量节点7传递过来的值
wire [5:0] value_check_8_to_variable_7;
wire enable_check_8_to_variable_7;
wire [5:0] value_variable_7_to_check_8;
wire enable_variable_7_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_7 = value_check_8_to_variable[5:0];
assign enable_check_8_to_variable_7 = enable_check_8_to_variable[0];
// 对变量节点7传递过来的值进行组合
assign value_variable_to_check_8[5:0] = value_variable_7_to_check_8;
assign enable_variable_to_check_8[0] = enable_variable_7_to_check_8;

// 拆分后校验节点8传递给变量节点49的值以及对变量节点49传递过来的值
wire [5:0] value_check_8_to_variable_49;
wire enable_check_8_to_variable_49;
wire [5:0] value_variable_49_to_check_8;
wire enable_variable_49_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_49 = value_check_8_to_variable[11:6];
assign enable_check_8_to_variable_49 = enable_check_8_to_variable[1];
// 对变量节点49传递过来的值进行组合
assign value_variable_to_check_8[11:6] = value_variable_49_to_check_8;
assign enable_variable_to_check_8[1] = enable_variable_49_to_check_8;

// 拆分后校验节点8传递给变量节点94的值以及对变量节点94传递过来的值
wire [5:0] value_check_8_to_variable_94;
wire enable_check_8_to_variable_94;
wire [5:0] value_variable_94_to_check_8;
wire enable_variable_94_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_94 = value_check_8_to_variable[17:12];
assign enable_check_8_to_variable_94 = enable_check_8_to_variable[2];
// 对变量节点94传递过来的值进行组合
assign value_variable_to_check_8[17:12] = value_variable_94_to_check_8;
assign enable_variable_to_check_8[2] = enable_variable_94_to_check_8;

// 拆分后校验节点8传递给变量节点137的值以及对变量节点137传递过来的值
wire [5:0] value_check_8_to_variable_137;
wire enable_check_8_to_variable_137;
wire [5:0] value_variable_137_to_check_8;
wire enable_variable_137_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_137 = value_check_8_to_variable[23:18];
assign enable_check_8_to_variable_137 = enable_check_8_to_variable[3];
// 对变量节点137传递过来的值进行组合
assign value_variable_to_check_8[23:18] = value_variable_137_to_check_8;
assign enable_variable_to_check_8[3] = enable_variable_137_to_check_8;

// 拆分后校验节点8传递给变量节点180的值以及对变量节点180传递过来的值
wire [5:0] value_check_8_to_variable_180;
wire enable_check_8_to_variable_180;
wire [5:0] value_variable_180_to_check_8;
wire enable_variable_180_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_180 = value_check_8_to_variable[29:24];
assign enable_check_8_to_variable_180 = enable_check_8_to_variable[4];
// 对变量节点180传递过来的值进行组合
assign value_variable_to_check_8[29:24] = value_variable_180_to_check_8;
assign enable_variable_to_check_8[4] = enable_variable_180_to_check_8;

// 拆分后校验节点8传递给变量节点222的值以及对变量节点222传递过来的值
wire [5:0] value_check_8_to_variable_222;
wire enable_check_8_to_variable_222;
wire [5:0] value_variable_222_to_check_8;
wire enable_variable_222_to_check_8;
// 对校验节点8的输出值进行拆分
assign value_check_8_to_variable_222 = value_check_8_to_variable[35:30];
assign enable_check_8_to_variable_222 = enable_check_8_to_variable[5];
// 对变量节点222传递过来的值进行组合
assign value_variable_to_check_8[35:30] = value_variable_222_to_check_8;
assign enable_variable_to_check_8[5] = enable_variable_222_to_check_8;


// 校验节点9的接口
wire [35:0] value_variable_to_check_9;
wire [35:0] value_check_9_to_variable;
wire [5:0] enable_variable_to_check_9;
wire [5:0] enable_check_9_to_variable;

// 拆分后校验节点9传递给变量节点8的值以及对变量节点8传递过来的值
wire [5:0] value_check_9_to_variable_8;
wire enable_check_9_to_variable_8;
wire [5:0] value_variable_8_to_check_9;
wire enable_variable_8_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_8 = value_check_9_to_variable[5:0];
assign enable_check_9_to_variable_8 = enable_check_9_to_variable[0];
// 对变量节点8传递过来的值进行组合
assign value_variable_to_check_9[5:0] = value_variable_8_to_check_9;
assign enable_variable_to_check_9[0] = enable_variable_8_to_check_9;

// 拆分后校验节点9传递给变量节点50的值以及对变量节点50传递过来的值
wire [5:0] value_check_9_to_variable_50;
wire enable_check_9_to_variable_50;
wire [5:0] value_variable_50_to_check_9;
wire enable_variable_50_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_50 = value_check_9_to_variable[11:6];
assign enable_check_9_to_variable_50 = enable_check_9_to_variable[1];
// 对变量节点50传递过来的值进行组合
assign value_variable_to_check_9[11:6] = value_variable_50_to_check_9;
assign enable_variable_to_check_9[1] = enable_variable_50_to_check_9;

// 拆分后校验节点9传递给变量节点95的值以及对变量节点95传递过来的值
wire [5:0] value_check_9_to_variable_95;
wire enable_check_9_to_variable_95;
wire [5:0] value_variable_95_to_check_9;
wire enable_variable_95_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_95 = value_check_9_to_variable[17:12];
assign enable_check_9_to_variable_95 = enable_check_9_to_variable[2];
// 对变量节点95传递过来的值进行组合
assign value_variable_to_check_9[17:12] = value_variable_95_to_check_9;
assign enable_variable_to_check_9[2] = enable_variable_95_to_check_9;

// 拆分后校验节点9传递给变量节点138的值以及对变量节点138传递过来的值
wire [5:0] value_check_9_to_variable_138;
wire enable_check_9_to_variable_138;
wire [5:0] value_variable_138_to_check_9;
wire enable_variable_138_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_138 = value_check_9_to_variable[23:18];
assign enable_check_9_to_variable_138 = enable_check_9_to_variable[3];
// 对变量节点138传递过来的值进行组合
assign value_variable_to_check_9[23:18] = value_variable_138_to_check_9;
assign enable_variable_to_check_9[3] = enable_variable_138_to_check_9;

// 拆分后校验节点9传递给变量节点179的值以及对变量节点179传递过来的值
wire [5:0] value_check_9_to_variable_179;
wire enable_check_9_to_variable_179;
wire [5:0] value_variable_179_to_check_9;
wire enable_variable_179_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_179 = value_check_9_to_variable[29:24];
assign enable_check_9_to_variable_179 = enable_check_9_to_variable[4];
// 对变量节点179传递过来的值进行组合
assign value_variable_to_check_9[29:24] = value_variable_179_to_check_9;
assign enable_variable_to_check_9[4] = enable_variable_179_to_check_9;

// 拆分后校验节点9传递给变量节点223的值以及对变量节点223传递过来的值
wire [5:0] value_check_9_to_variable_223;
wire enable_check_9_to_variable_223;
wire [5:0] value_variable_223_to_check_9;
wire enable_variable_223_to_check_9;
// 对校验节点9的输出值进行拆分
assign value_check_9_to_variable_223 = value_check_9_to_variable[35:30];
assign enable_check_9_to_variable_223 = enable_check_9_to_variable[5];
// 对变量节点223传递过来的值进行组合
assign value_variable_to_check_9[35:30] = value_variable_223_to_check_9;
assign enable_variable_to_check_9[5] = enable_variable_223_to_check_9;


// 校验节点10的接口
wire [35:0] value_variable_to_check_10;
wire [35:0] value_check_10_to_variable;
wire [5:0] enable_variable_to_check_10;
wire [5:0] enable_check_10_to_variable;

// 拆分后校验节点10传递给变量节点9的值以及对变量节点9传递过来的值
wire [5:0] value_check_10_to_variable_9;
wire enable_check_10_to_variable_9;
wire [5:0] value_variable_9_to_check_10;
wire enable_variable_9_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_9 = value_check_10_to_variable[5:0];
assign enable_check_10_to_variable_9 = enable_check_10_to_variable[0];
// 对变量节点9传递过来的值进行组合
assign value_variable_to_check_10[5:0] = value_variable_9_to_check_10;
assign enable_variable_to_check_10[0] = enable_variable_9_to_check_10;

// 拆分后校验节点10传递给变量节点51的值以及对变量节点51传递过来的值
wire [5:0] value_check_10_to_variable_51;
wire enable_check_10_to_variable_51;
wire [5:0] value_variable_51_to_check_10;
wire enable_variable_51_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_51 = value_check_10_to_variable[11:6];
assign enable_check_10_to_variable_51 = enable_check_10_to_variable[1];
// 对变量节点51传递过来的值进行组合
assign value_variable_to_check_10[11:6] = value_variable_51_to_check_10;
assign enable_variable_to_check_10[1] = enable_variable_51_to_check_10;

// 拆分后校验节点10传递给变量节点96的值以及对变量节点96传递过来的值
wire [5:0] value_check_10_to_variable_96;
wire enable_check_10_to_variable_96;
wire [5:0] value_variable_96_to_check_10;
wire enable_variable_96_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_96 = value_check_10_to_variable[17:12];
assign enable_check_10_to_variable_96 = enable_check_10_to_variable[2];
// 对变量节点96传递过来的值进行组合
assign value_variable_to_check_10[17:12] = value_variable_96_to_check_10;
assign enable_variable_to_check_10[2] = enable_variable_96_to_check_10;

// 拆分后校验节点10传递给变量节点139的值以及对变量节点139传递过来的值
wire [5:0] value_check_10_to_variable_139;
wire enable_check_10_to_variable_139;
wire [5:0] value_variable_139_to_check_10;
wire enable_variable_139_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_139 = value_check_10_to_variable[23:18];
assign enable_check_10_to_variable_139 = enable_check_10_to_variable[3];
// 对变量节点139传递过来的值进行组合
assign value_variable_to_check_10[23:18] = value_variable_139_to_check_10;
assign enable_variable_to_check_10[3] = enable_variable_139_to_check_10;

// 拆分后校验节点10传递给变量节点181的值以及对变量节点181传递过来的值
wire [5:0] value_check_10_to_variable_181;
wire enable_check_10_to_variable_181;
wire [5:0] value_variable_181_to_check_10;
wire enable_variable_181_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_181 = value_check_10_to_variable[29:24];
assign enable_check_10_to_variable_181 = enable_check_10_to_variable[4];
// 对变量节点181传递过来的值进行组合
assign value_variable_to_check_10[29:24] = value_variable_181_to_check_10;
assign enable_variable_to_check_10[4] = enable_variable_181_to_check_10;

// 拆分后校验节点10传递给变量节点222的值以及对变量节点222传递过来的值
wire [5:0] value_check_10_to_variable_222;
wire enable_check_10_to_variable_222;
wire [5:0] value_variable_222_to_check_10;
wire enable_variable_222_to_check_10;
// 对校验节点10的输出值进行拆分
assign value_check_10_to_variable_222 = value_check_10_to_variable[35:30];
assign enable_check_10_to_variable_222 = enable_check_10_to_variable[5];
// 对变量节点222传递过来的值进行组合
assign value_variable_to_check_10[35:30] = value_variable_222_to_check_10;
assign enable_variable_to_check_10[5] = enable_variable_222_to_check_10;


// 校验节点11的接口
wire [35:0] value_variable_to_check_11;
wire [35:0] value_check_11_to_variable;
wire [5:0] enable_variable_to_check_11;
wire [5:0] enable_check_11_to_variable;

// 拆分后校验节点11传递给变量节点10的值以及对变量节点10传递过来的值
wire [5:0] value_check_11_to_variable_10;
wire enable_check_11_to_variable_10;
wire [5:0] value_variable_10_to_check_11;
wire enable_variable_10_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_10 = value_check_11_to_variable[5:0];
assign enable_check_11_to_variable_10 = enable_check_11_to_variable[0];
// 对变量节点10传递过来的值进行组合
assign value_variable_to_check_11[5:0] = value_variable_10_to_check_11;
assign enable_variable_to_check_11[0] = enable_variable_10_to_check_11;

// 拆分后校验节点11传递给变量节点52的值以及对变量节点52传递过来的值
wire [5:0] value_check_11_to_variable_52;
wire enable_check_11_to_variable_52;
wire [5:0] value_variable_52_to_check_11;
wire enable_variable_52_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_52 = value_check_11_to_variable[11:6];
assign enable_check_11_to_variable_52 = enable_check_11_to_variable[1];
// 对变量节点52传递过来的值进行组合
assign value_variable_to_check_11[11:6] = value_variable_52_to_check_11;
assign enable_variable_to_check_11[1] = enable_variable_52_to_check_11;

// 拆分后校验节点11传递给变量节点97的值以及对变量节点97传递过来的值
wire [5:0] value_check_11_to_variable_97;
wire enable_check_11_to_variable_97;
wire [5:0] value_variable_97_to_check_11;
wire enable_variable_97_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_97 = value_check_11_to_variable[17:12];
assign enable_check_11_to_variable_97 = enable_check_11_to_variable[2];
// 对变量节点97传递过来的值进行组合
assign value_variable_to_check_11[17:12] = value_variable_97_to_check_11;
assign enable_variable_to_check_11[2] = enable_variable_97_to_check_11;

// 拆分后校验节点11传递给变量节点140的值以及对变量节点140传递过来的值
wire [5:0] value_check_11_to_variable_140;
wire enable_check_11_to_variable_140;
wire [5:0] value_variable_140_to_check_11;
wire enable_variable_140_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_140 = value_check_11_to_variable[23:18];
assign enable_check_11_to_variable_140 = enable_check_11_to_variable[3];
// 对变量节点140传递过来的值进行组合
assign value_variable_to_check_11[23:18] = value_variable_140_to_check_11;
assign enable_variable_to_check_11[3] = enable_variable_140_to_check_11;

// 拆分后校验节点11传递给变量节点182的值以及对变量节点182传递过来的值
wire [5:0] value_check_11_to_variable_182;
wire enable_check_11_to_variable_182;
wire [5:0] value_variable_182_to_check_11;
wire enable_variable_182_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_182 = value_check_11_to_variable[29:24];
assign enable_check_11_to_variable_182 = enable_check_11_to_variable[4];
// 对变量节点182传递过来的值进行组合
assign value_variable_to_check_11[29:24] = value_variable_182_to_check_11;
assign enable_variable_to_check_11[4] = enable_variable_182_to_check_11;

// 拆分后校验节点11传递给变量节点224的值以及对变量节点224传递过来的值
wire [5:0] value_check_11_to_variable_224;
wire enable_check_11_to_variable_224;
wire [5:0] value_variable_224_to_check_11;
wire enable_variable_224_to_check_11;
// 对校验节点11的输出值进行拆分
assign value_check_11_to_variable_224 = value_check_11_to_variable[35:30];
assign enable_check_11_to_variable_224 = enable_check_11_to_variable[5];
// 对变量节点224传递过来的值进行组合
assign value_variable_to_check_11[35:30] = value_variable_224_to_check_11;
assign enable_variable_to_check_11[5] = enable_variable_224_to_check_11;


// 校验节点12的接口
wire [35:0] value_variable_to_check_12;
wire [35:0] value_check_12_to_variable;
wire [5:0] enable_variable_to_check_12;
wire [5:0] enable_check_12_to_variable;

// 拆分后校验节点12传递给变量节点11的值以及对变量节点11传递过来的值
wire [5:0] value_check_12_to_variable_11;
wire enable_check_12_to_variable_11;
wire [5:0] value_variable_11_to_check_12;
wire enable_variable_11_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_11 = value_check_12_to_variable[5:0];
assign enable_check_12_to_variable_11 = enable_check_12_to_variable[0];
// 对变量节点11传递过来的值进行组合
assign value_variable_to_check_12[5:0] = value_variable_11_to_check_12;
assign enable_variable_to_check_12[0] = enable_variable_11_to_check_12;

// 拆分后校验节点12传递给变量节点53的值以及对变量节点53传递过来的值
wire [5:0] value_check_12_to_variable_53;
wire enable_check_12_to_variable_53;
wire [5:0] value_variable_53_to_check_12;
wire enable_variable_53_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_53 = value_check_12_to_variable[11:6];
assign enable_check_12_to_variable_53 = enable_check_12_to_variable[1];
// 对变量节点53传递过来的值进行组合
assign value_variable_to_check_12[11:6] = value_variable_53_to_check_12;
assign enable_variable_to_check_12[1] = enable_variable_53_to_check_12;

// 拆分后校验节点12传递给变量节点98的值以及对变量节点98传递过来的值
wire [5:0] value_check_12_to_variable_98;
wire enable_check_12_to_variable_98;
wire [5:0] value_variable_98_to_check_12;
wire enable_variable_98_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_98 = value_check_12_to_variable[17:12];
assign enable_check_12_to_variable_98 = enable_check_12_to_variable[2];
// 对变量节点98传递过来的值进行组合
assign value_variable_to_check_12[17:12] = value_variable_98_to_check_12;
assign enable_variable_to_check_12[2] = enable_variable_98_to_check_12;

// 拆分后校验节点12传递给变量节点112的值以及对变量节点112传递过来的值
wire [5:0] value_check_12_to_variable_112;
wire enable_check_12_to_variable_112;
wire [5:0] value_variable_112_to_check_12;
wire enable_variable_112_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_112 = value_check_12_to_variable[23:18];
assign enable_check_12_to_variable_112 = enable_check_12_to_variable[3];
// 对变量节点112传递过来的值进行组合
assign value_variable_to_check_12[23:18] = value_variable_112_to_check_12;
assign enable_variable_to_check_12[3] = enable_variable_112_to_check_12;

// 拆分后校验节点12传递给变量节点183的值以及对变量节点183传递过来的值
wire [5:0] value_check_12_to_variable_183;
wire enable_check_12_to_variable_183;
wire [5:0] value_variable_183_to_check_12;
wire enable_variable_183_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_183 = value_check_12_to_variable[29:24];
assign enable_check_12_to_variable_183 = enable_check_12_to_variable[4];
// 对变量节点183传递过来的值进行组合
assign value_variable_to_check_12[29:24] = value_variable_183_to_check_12;
assign enable_variable_to_check_12[4] = enable_variable_183_to_check_12;

// 拆分后校验节点12传递给变量节点225的值以及对变量节点225传递过来的值
wire [5:0] value_check_12_to_variable_225;
wire enable_check_12_to_variable_225;
wire [5:0] value_variable_225_to_check_12;
wire enable_variable_225_to_check_12;
// 对校验节点12的输出值进行拆分
assign value_check_12_to_variable_225 = value_check_12_to_variable[35:30];
assign enable_check_12_to_variable_225 = enable_check_12_to_variable[5];
// 对变量节点225传递过来的值进行组合
assign value_variable_to_check_12[35:30] = value_variable_225_to_check_12;
assign enable_variable_to_check_12[5] = enable_variable_225_to_check_12;


// 校验节点13的接口
wire [35:0] value_variable_to_check_13;
wire [35:0] value_check_13_to_variable;
wire [5:0] enable_variable_to_check_13;
wire [5:0] enable_check_13_to_variable;

// 拆分后校验节点13传递给变量节点12的值以及对变量节点12传递过来的值
wire [5:0] value_check_13_to_variable_12;
wire enable_check_13_to_variable_12;
wire [5:0] value_variable_12_to_check_13;
wire enable_variable_12_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_12 = value_check_13_to_variable[5:0];
assign enable_check_13_to_variable_12 = enable_check_13_to_variable[0];
// 对变量节点12传递过来的值进行组合
assign value_variable_to_check_13[5:0] = value_variable_12_to_check_13;
assign enable_variable_to_check_13[0] = enable_variable_12_to_check_13;

// 拆分后校验节点13传递给变量节点54的值以及对变量节点54传递过来的值
wire [5:0] value_check_13_to_variable_54;
wire enable_check_13_to_variable_54;
wire [5:0] value_variable_54_to_check_13;
wire enable_variable_54_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_54 = value_check_13_to_variable[11:6];
assign enable_check_13_to_variable_54 = enable_check_13_to_variable[1];
// 对变量节点54传递过来的值进行组合
assign value_variable_to_check_13[11:6] = value_variable_54_to_check_13;
assign enable_variable_to_check_13[1] = enable_variable_54_to_check_13;

// 拆分后校验节点13传递给变量节点99的值以及对变量节点99传递过来的值
wire [5:0] value_check_13_to_variable_99;
wire enable_check_13_to_variable_99;
wire [5:0] value_variable_99_to_check_13;
wire enable_variable_99_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_99 = value_check_13_to_variable[17:12];
assign enable_check_13_to_variable_99 = enable_check_13_to_variable[2];
// 对变量节点99传递过来的值进行组合
assign value_variable_to_check_13[17:12] = value_variable_99_to_check_13;
assign enable_variable_to_check_13[2] = enable_variable_99_to_check_13;

// 拆分后校验节点13传递给变量节点141的值以及对变量节点141传递过来的值
wire [5:0] value_check_13_to_variable_141;
wire enable_check_13_to_variable_141;
wire [5:0] value_variable_141_to_check_13;
wire enable_variable_141_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_141 = value_check_13_to_variable[23:18];
assign enable_check_13_to_variable_141 = enable_check_13_to_variable[3];
// 对变量节点141传递过来的值进行组合
assign value_variable_to_check_13[23:18] = value_variable_141_to_check_13;
assign enable_variable_to_check_13[3] = enable_variable_141_to_check_13;

// 拆分后校验节点13传递给变量节点184的值以及对变量节点184传递过来的值
wire [5:0] value_check_13_to_variable_184;
wire enable_check_13_to_variable_184;
wire [5:0] value_variable_184_to_check_13;
wire enable_variable_184_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_184 = value_check_13_to_variable[29:24];
assign enable_check_13_to_variable_184 = enable_check_13_to_variable[4];
// 对变量节点184传递过来的值进行组合
assign value_variable_to_check_13[29:24] = value_variable_184_to_check_13;
assign enable_variable_to_check_13[4] = enable_variable_184_to_check_13;

// 拆分后校验节点13传递给变量节点226的值以及对变量节点226传递过来的值
wire [5:0] value_check_13_to_variable_226;
wire enable_check_13_to_variable_226;
wire [5:0] value_variable_226_to_check_13;
wire enable_variable_226_to_check_13;
// 对校验节点13的输出值进行拆分
assign value_check_13_to_variable_226 = value_check_13_to_variable[35:30];
assign enable_check_13_to_variable_226 = enable_check_13_to_variable[5];
// 对变量节点226传递过来的值进行组合
assign value_variable_to_check_13[35:30] = value_variable_226_to_check_13;
assign enable_variable_to_check_13[5] = enable_variable_226_to_check_13;


// 校验节点14的接口
wire [35:0] value_variable_to_check_14;
wire [35:0] value_check_14_to_variable;
wire [5:0] enable_variable_to_check_14;
wire [5:0] enable_check_14_to_variable;

// 拆分后校验节点14传递给变量节点9的值以及对变量节点9传递过来的值
wire [5:0] value_check_14_to_variable_9;
wire enable_check_14_to_variable_9;
wire [5:0] value_variable_9_to_check_14;
wire enable_variable_9_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_9 = value_check_14_to_variable[5:0];
assign enable_check_14_to_variable_9 = enable_check_14_to_variable[0];
// 对变量节点9传递过来的值进行组合
assign value_variable_to_check_14[5:0] = value_variable_9_to_check_14;
assign enable_variable_to_check_14[0] = enable_variable_9_to_check_14;

// 拆分后校验节点14传递给变量节点55的值以及对变量节点55传递过来的值
wire [5:0] value_check_14_to_variable_55;
wire enable_check_14_to_variable_55;
wire [5:0] value_variable_55_to_check_14;
wire enable_variable_55_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_55 = value_check_14_to_variable[11:6];
assign enable_check_14_to_variable_55 = enable_check_14_to_variable[1];
// 对变量节点55传递过来的值进行组合
assign value_variable_to_check_14[11:6] = value_variable_55_to_check_14;
assign enable_variable_to_check_14[1] = enable_variable_55_to_check_14;

// 拆分后校验节点14传递给变量节点100的值以及对变量节点100传递过来的值
wire [5:0] value_check_14_to_variable_100;
wire enable_check_14_to_variable_100;
wire [5:0] value_variable_100_to_check_14;
wire enable_variable_100_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_100 = value_check_14_to_variable[17:12];
assign enable_check_14_to_variable_100 = enable_check_14_to_variable[2];
// 对变量节点100传递过来的值进行组合
assign value_variable_to_check_14[17:12] = value_variable_100_to_check_14;
assign enable_variable_to_check_14[2] = enable_variable_100_to_check_14;

// 拆分后校验节点14传递给变量节点142的值以及对变量节点142传递过来的值
wire [5:0] value_check_14_to_variable_142;
wire enable_check_14_to_variable_142;
wire [5:0] value_variable_142_to_check_14;
wire enable_variable_142_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_142 = value_check_14_to_variable[23:18];
assign enable_check_14_to_variable_142 = enable_check_14_to_variable[3];
// 对变量节点142传递过来的值进行组合
assign value_variable_to_check_14[23:18] = value_variable_142_to_check_14;
assign enable_variable_to_check_14[3] = enable_variable_142_to_check_14;

// 拆分后校验节点14传递给变量节点185的值以及对变量节点185传递过来的值
wire [5:0] value_check_14_to_variable_185;
wire enable_check_14_to_variable_185;
wire [5:0] value_variable_185_to_check_14;
wire enable_variable_185_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_185 = value_check_14_to_variable[29:24];
assign enable_check_14_to_variable_185 = enable_check_14_to_variable[4];
// 对变量节点185传递过来的值进行组合
assign value_variable_to_check_14[29:24] = value_variable_185_to_check_14;
assign enable_variable_to_check_14[4] = enable_variable_185_to_check_14;

// 拆分后校验节点14传递给变量节点227的值以及对变量节点227传递过来的值
wire [5:0] value_check_14_to_variable_227;
wire enable_check_14_to_variable_227;
wire [5:0] value_variable_227_to_check_14;
wire enable_variable_227_to_check_14;
// 对校验节点14的输出值进行拆分
assign value_check_14_to_variable_227 = value_check_14_to_variable[35:30];
assign enable_check_14_to_variable_227 = enable_check_14_to_variable[5];
// 对变量节点227传递过来的值进行组合
assign value_variable_to_check_14[35:30] = value_variable_227_to_check_14;
assign enable_variable_to_check_14[5] = enable_variable_227_to_check_14;


// 校验节点15的接口
wire [35:0] value_variable_to_check_15;
wire [35:0] value_check_15_to_variable;
wire [5:0] enable_variable_to_check_15;
wire [5:0] enable_check_15_to_variable;

// 拆分后校验节点15传递给变量节点12的值以及对变量节点12传递过来的值
wire [5:0] value_check_15_to_variable_12;
wire enable_check_15_to_variable_12;
wire [5:0] value_variable_12_to_check_15;
wire enable_variable_12_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_12 = value_check_15_to_variable[5:0];
assign enable_check_15_to_variable_12 = enable_check_15_to_variable[0];
// 对变量节点12传递过来的值进行组合
assign value_variable_to_check_15[5:0] = value_variable_12_to_check_15;
assign enable_variable_to_check_15[0] = enable_variable_12_to_check_15;

// 拆分后校验节点15传递给变量节点56的值以及对变量节点56传递过来的值
wire [5:0] value_check_15_to_variable_56;
wire enable_check_15_to_variable_56;
wire [5:0] value_variable_56_to_check_15;
wire enable_variable_56_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_56 = value_check_15_to_variable[11:6];
assign enable_check_15_to_variable_56 = enable_check_15_to_variable[1];
// 对变量节点56传递过来的值进行组合
assign value_variable_to_check_15[11:6] = value_variable_56_to_check_15;
assign enable_variable_to_check_15[1] = enable_variable_56_to_check_15;

// 拆分后校验节点15传递给变量节点101的值以及对变量节点101传递过来的值
wire [5:0] value_check_15_to_variable_101;
wire enable_check_15_to_variable_101;
wire [5:0] value_variable_101_to_check_15;
wire enable_variable_101_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_101 = value_check_15_to_variable[17:12];
assign enable_check_15_to_variable_101 = enable_check_15_to_variable[2];
// 对变量节点101传递过来的值进行组合
assign value_variable_to_check_15[17:12] = value_variable_101_to_check_15;
assign enable_variable_to_check_15[2] = enable_variable_101_to_check_15;

// 拆分后校验节点15传递给变量节点143的值以及对变量节点143传递过来的值
wire [5:0] value_check_15_to_variable_143;
wire enable_check_15_to_variable_143;
wire [5:0] value_variable_143_to_check_15;
wire enable_variable_143_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_143 = value_check_15_to_variable[23:18];
assign enable_check_15_to_variable_143 = enable_check_15_to_variable[3];
// 对变量节点143传递过来的值进行组合
assign value_variable_to_check_15[23:18] = value_variable_143_to_check_15;
assign enable_variable_to_check_15[3] = enable_variable_143_to_check_15;

// 拆分后校验节点15传递给变量节点186的值以及对变量节点186传递过来的值
wire [5:0] value_check_15_to_variable_186;
wire enable_check_15_to_variable_186;
wire [5:0] value_variable_186_to_check_15;
wire enable_variable_186_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_186 = value_check_15_to_variable[29:24];
assign enable_check_15_to_variable_186 = enable_check_15_to_variable[4];
// 对变量节点186传递过来的值进行组合
assign value_variable_to_check_15[29:24] = value_variable_186_to_check_15;
assign enable_variable_to_check_15[4] = enable_variable_186_to_check_15;

// 拆分后校验节点15传递给变量节点217的值以及对变量节点217传递过来的值
wire [5:0] value_check_15_to_variable_217;
wire enable_check_15_to_variable_217;
wire [5:0] value_variable_217_to_check_15;
wire enable_variable_217_to_check_15;
// 对校验节点15的输出值进行拆分
assign value_check_15_to_variable_217 = value_check_15_to_variable[35:30];
assign enable_check_15_to_variable_217 = enable_check_15_to_variable[5];
// 对变量节点217传递过来的值进行组合
assign value_variable_to_check_15[35:30] = value_variable_217_to_check_15;
assign enable_variable_to_check_15[5] = enable_variable_217_to_check_15;


// 校验节点16的接口
wire [35:0] value_variable_to_check_16;
wire [35:0] value_check_16_to_variable;
wire [5:0] enable_variable_to_check_16;
wire [5:0] enable_check_16_to_variable;

// 拆分后校验节点16传递给变量节点13的值以及对变量节点13传递过来的值
wire [5:0] value_check_16_to_variable_13;
wire enable_check_16_to_variable_13;
wire [5:0] value_variable_13_to_check_16;
wire enable_variable_13_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_13 = value_check_16_to_variable[5:0];
assign enable_check_16_to_variable_13 = enable_check_16_to_variable[0];
// 对变量节点13传递过来的值进行组合
assign value_variable_to_check_16[5:0] = value_variable_13_to_check_16;
assign enable_variable_to_check_16[0] = enable_variable_13_to_check_16;

// 拆分后校验节点16传递给变量节点57的值以及对变量节点57传递过来的值
wire [5:0] value_check_16_to_variable_57;
wire enable_check_16_to_variable_57;
wire [5:0] value_variable_57_to_check_16;
wire enable_variable_57_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_57 = value_check_16_to_variable[11:6];
assign enable_check_16_to_variable_57 = enable_check_16_to_variable[1];
// 对变量节点57传递过来的值进行组合
assign value_variable_to_check_16[11:6] = value_variable_57_to_check_16;
assign enable_variable_to_check_16[1] = enable_variable_57_to_check_16;

// 拆分后校验节点16传递给变量节点102的值以及对变量节点102传递过来的值
wire [5:0] value_check_16_to_variable_102;
wire enable_check_16_to_variable_102;
wire [5:0] value_variable_102_to_check_16;
wire enable_variable_102_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_102 = value_check_16_to_variable[17:12];
assign enable_check_16_to_variable_102 = enable_check_16_to_variable[2];
// 对变量节点102传递过来的值进行组合
assign value_variable_to_check_16[17:12] = value_variable_102_to_check_16;
assign enable_variable_to_check_16[2] = enable_variable_102_to_check_16;

// 拆分后校验节点16传递给变量节点144的值以及对变量节点144传递过来的值
wire [5:0] value_check_16_to_variable_144;
wire enable_check_16_to_variable_144;
wire [5:0] value_variable_144_to_check_16;
wire enable_variable_144_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_144 = value_check_16_to_variable[23:18];
assign enable_check_16_to_variable_144 = enable_check_16_to_variable[3];
// 对变量节点144传递过来的值进行组合
assign value_variable_to_check_16[23:18] = value_variable_144_to_check_16;
assign enable_variable_to_check_16[3] = enable_variable_144_to_check_16;

// 拆分后校验节点16传递给变量节点184的值以及对变量节点184传递过来的值
wire [5:0] value_check_16_to_variable_184;
wire enable_check_16_to_variable_184;
wire [5:0] value_variable_184_to_check_16;
wire enable_variable_184_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_184 = value_check_16_to_variable[29:24];
assign enable_check_16_to_variable_184 = enable_check_16_to_variable[4];
// 对变量节点184传递过来的值进行组合
assign value_variable_to_check_16[29:24] = value_variable_184_to_check_16;
assign enable_variable_to_check_16[4] = enable_variable_184_to_check_16;

// 拆分后校验节点16传递给变量节点216的值以及对变量节点216传递过来的值
wire [5:0] value_check_16_to_variable_216;
wire enable_check_16_to_variable_216;
wire [5:0] value_variable_216_to_check_16;
wire enable_variable_216_to_check_16;
// 对校验节点16的输出值进行拆分
assign value_check_16_to_variable_216 = value_check_16_to_variable[35:30];
assign enable_check_16_to_variable_216 = enable_check_16_to_variable[5];
// 对变量节点216传递过来的值进行组合
assign value_variable_to_check_16[35:30] = value_variable_216_to_check_16;
assign enable_variable_to_check_16[5] = enable_variable_216_to_check_16;


// 校验节点17的接口
wire [35:0] value_variable_to_check_17;
wire [35:0] value_check_17_to_variable;
wire [5:0] enable_variable_to_check_17;
wire [5:0] enable_check_17_to_variable;

// 拆分后校验节点17传递给变量节点14的值以及对变量节点14传递过来的值
wire [5:0] value_check_17_to_variable_14;
wire enable_check_17_to_variable_14;
wire [5:0] value_variable_14_to_check_17;
wire enable_variable_14_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_14 = value_check_17_to_variable[5:0];
assign enable_check_17_to_variable_14 = enable_check_17_to_variable[0];
// 对变量节点14传递过来的值进行组合
assign value_variable_to_check_17[5:0] = value_variable_14_to_check_17;
assign enable_variable_to_check_17[0] = enable_variable_14_to_check_17;

// 拆分后校验节点17传递给变量节点58的值以及对变量节点58传递过来的值
wire [5:0] value_check_17_to_variable_58;
wire enable_check_17_to_variable_58;
wire [5:0] value_variable_58_to_check_17;
wire enable_variable_58_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_58 = value_check_17_to_variable[11:6];
assign enable_check_17_to_variable_58 = enable_check_17_to_variable[1];
// 对变量节点58传递过来的值进行组合
assign value_variable_to_check_17[11:6] = value_variable_58_to_check_17;
assign enable_variable_to_check_17[1] = enable_variable_58_to_check_17;

// 拆分后校验节点17传递给变量节点102的值以及对变量节点102传递过来的值
wire [5:0] value_check_17_to_variable_102;
wire enable_check_17_to_variable_102;
wire [5:0] value_variable_102_to_check_17;
wire enable_variable_102_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_102 = value_check_17_to_variable[17:12];
assign enable_check_17_to_variable_102 = enable_check_17_to_variable[2];
// 对变量节点102传递过来的值进行组合
assign value_variable_to_check_17[17:12] = value_variable_102_to_check_17;
assign enable_variable_to_check_17[2] = enable_variable_102_to_check_17;

// 拆分后校验节点17传递给变量节点145的值以及对变量节点145传递过来的值
wire [5:0] value_check_17_to_variable_145;
wire enable_check_17_to_variable_145;
wire [5:0] value_variable_145_to_check_17;
wire enable_variable_145_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_145 = value_check_17_to_variable[23:18];
assign enable_check_17_to_variable_145 = enable_check_17_to_variable[3];
// 对变量节点145传递过来的值进行组合
assign value_variable_to_check_17[23:18] = value_variable_145_to_check_17;
assign enable_variable_to_check_17[3] = enable_variable_145_to_check_17;

// 拆分后校验节点17传递给变量节点187的值以及对变量节点187传递过来的值
wire [5:0] value_check_17_to_variable_187;
wire enable_check_17_to_variable_187;
wire [5:0] value_variable_187_to_check_17;
wire enable_variable_187_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_187 = value_check_17_to_variable[29:24];
assign enable_check_17_to_variable_187 = enable_check_17_to_variable[4];
// 对变量节点187传递过来的值进行组合
assign value_variable_to_check_17[29:24] = value_variable_187_to_check_17;
assign enable_variable_to_check_17[4] = enable_variable_187_to_check_17;

// 拆分后校验节点17传递给变量节点228的值以及对变量节点228传递过来的值
wire [5:0] value_check_17_to_variable_228;
wire enable_check_17_to_variable_228;
wire [5:0] value_variable_228_to_check_17;
wire enable_variable_228_to_check_17;
// 对校验节点17的输出值进行拆分
assign value_check_17_to_variable_228 = value_check_17_to_variable[35:30];
assign enable_check_17_to_variable_228 = enable_check_17_to_variable[5];
// 对变量节点228传递过来的值进行组合
assign value_variable_to_check_17[35:30] = value_variable_228_to_check_17;
assign enable_variable_to_check_17[5] = enable_variable_228_to_check_17;


// 校验节点18的接口
wire [35:0] value_variable_to_check_18;
wire [35:0] value_check_18_to_variable;
wire [5:0] enable_variable_to_check_18;
wire [5:0] enable_check_18_to_variable;

// 拆分后校验节点18传递给变量节点15的值以及对变量节点15传递过来的值
wire [5:0] value_check_18_to_variable_15;
wire enable_check_18_to_variable_15;
wire [5:0] value_variable_15_to_check_18;
wire enable_variable_15_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_15 = value_check_18_to_variable[5:0];
assign enable_check_18_to_variable_15 = enable_check_18_to_variable[0];
// 对变量节点15传递过来的值进行组合
assign value_variable_to_check_18[5:0] = value_variable_15_to_check_18;
assign enable_variable_to_check_18[0] = enable_variable_15_to_check_18;

// 拆分后校验节点18传递给变量节点59的值以及对变量节点59传递过来的值
wire [5:0] value_check_18_to_variable_59;
wire enable_check_18_to_variable_59;
wire [5:0] value_variable_59_to_check_18;
wire enable_variable_59_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_59 = value_check_18_to_variable[11:6];
assign enable_check_18_to_variable_59 = enable_check_18_to_variable[1];
// 对变量节点59传递过来的值进行组合
assign value_variable_to_check_18[11:6] = value_variable_59_to_check_18;
assign enable_variable_to_check_18[1] = enable_variable_59_to_check_18;

// 拆分后校验节点18传递给变量节点101的值以及对变量节点101传递过来的值
wire [5:0] value_check_18_to_variable_101;
wire enable_check_18_to_variable_101;
wire [5:0] value_variable_101_to_check_18;
wire enable_variable_101_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_101 = value_check_18_to_variable[17:12];
assign enable_check_18_to_variable_101 = enable_check_18_to_variable[2];
// 对变量节点101传递过来的值进行组合
assign value_variable_to_check_18[17:12] = value_variable_101_to_check_18;
assign enable_variable_to_check_18[2] = enable_variable_101_to_check_18;

// 拆分后校验节点18传递给变量节点145的值以及对变量节点145传递过来的值
wire [5:0] value_check_18_to_variable_145;
wire enable_check_18_to_variable_145;
wire [5:0] value_variable_145_to_check_18;
wire enable_variable_145_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_145 = value_check_18_to_variable[23:18];
assign enable_check_18_to_variable_145 = enable_check_18_to_variable[3];
// 对变量节点145传递过来的值进行组合
assign value_variable_to_check_18[23:18] = value_variable_145_to_check_18;
assign enable_variable_to_check_18[3] = enable_variable_145_to_check_18;

// 拆分后校验节点18传递给变量节点188的值以及对变量节点188传递过来的值
wire [5:0] value_check_18_to_variable_188;
wire enable_check_18_to_variable_188;
wire [5:0] value_variable_188_to_check_18;
wire enable_variable_188_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_188 = value_check_18_to_variable[29:24];
assign enable_check_18_to_variable_188 = enable_check_18_to_variable[4];
// 对变量节点188传递过来的值进行组合
assign value_variable_to_check_18[29:24] = value_variable_188_to_check_18;
assign enable_variable_to_check_18[4] = enable_variable_188_to_check_18;

// 拆分后校验节点18传递给变量节点229的值以及对变量节点229传递过来的值
wire [5:0] value_check_18_to_variable_229;
wire enable_check_18_to_variable_229;
wire [5:0] value_variable_229_to_check_18;
wire enable_variable_229_to_check_18;
// 对校验节点18的输出值进行拆分
assign value_check_18_to_variable_229 = value_check_18_to_variable[35:30];
assign enable_check_18_to_variable_229 = enable_check_18_to_variable[5];
// 对变量节点229传递过来的值进行组合
assign value_variable_to_check_18[35:30] = value_variable_229_to_check_18;
assign enable_variable_to_check_18[5] = enable_variable_229_to_check_18;


// 校验节点19的接口
wire [35:0] value_variable_to_check_19;
wire [35:0] value_check_19_to_variable;
wire [5:0] enable_variable_to_check_19;
wire [5:0] enable_check_19_to_variable;

// 拆分后校验节点19传递给变量节点16的值以及对变量节点16传递过来的值
wire [5:0] value_check_19_to_variable_16;
wire enable_check_19_to_variable_16;
wire [5:0] value_variable_16_to_check_19;
wire enable_variable_16_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_16 = value_check_19_to_variable[5:0];
assign enable_check_19_to_variable_16 = enable_check_19_to_variable[0];
// 对变量节点16传递过来的值进行组合
assign value_variable_to_check_19[5:0] = value_variable_16_to_check_19;
assign enable_variable_to_check_19[0] = enable_variable_16_to_check_19;

// 拆分后校验节点19传递给变量节点60的值以及对变量节点60传递过来的值
wire [5:0] value_check_19_to_variable_60;
wire enable_check_19_to_variable_60;
wire [5:0] value_variable_60_to_check_19;
wire enable_variable_60_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_60 = value_check_19_to_variable[11:6];
assign enable_check_19_to_variable_60 = enable_check_19_to_variable[1];
// 对变量节点60传递过来的值进行组合
assign value_variable_to_check_19[11:6] = value_variable_60_to_check_19;
assign enable_variable_to_check_19[1] = enable_variable_60_to_check_19;

// 拆分后校验节点19传递给变量节点92的值以及对变量节点92传递过来的值
wire [5:0] value_check_19_to_variable_92;
wire enable_check_19_to_variable_92;
wire [5:0] value_variable_92_to_check_19;
wire enable_variable_92_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_92 = value_check_19_to_variable[17:12];
assign enable_check_19_to_variable_92 = enable_check_19_to_variable[2];
// 对变量节点92传递过来的值进行组合
assign value_variable_to_check_19[17:12] = value_variable_92_to_check_19;
assign enable_variable_to_check_19[2] = enable_variable_92_to_check_19;

// 拆分后校验节点19传递给变量节点146的值以及对变量节点146传递过来的值
wire [5:0] value_check_19_to_variable_146;
wire enable_check_19_to_variable_146;
wire [5:0] value_variable_146_to_check_19;
wire enable_variable_146_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_146 = value_check_19_to_variable[23:18];
assign enable_check_19_to_variable_146 = enable_check_19_to_variable[3];
// 对变量节点146传递过来的值进行组合
assign value_variable_to_check_19[23:18] = value_variable_146_to_check_19;
assign enable_variable_to_check_19[3] = enable_variable_146_to_check_19;

// 拆分后校验节点19传递给变量节点186的值以及对变量节点186传递过来的值
wire [5:0] value_check_19_to_variable_186;
wire enable_check_19_to_variable_186;
wire [5:0] value_variable_186_to_check_19;
wire enable_variable_186_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_186 = value_check_19_to_variable[29:24];
assign enable_check_19_to_variable_186 = enable_check_19_to_variable[4];
// 对变量节点186传递过来的值进行组合
assign value_variable_to_check_19[29:24] = value_variable_186_to_check_19;
assign enable_variable_to_check_19[4] = enable_variable_186_to_check_19;

// 拆分后校验节点19传递给变量节点230的值以及对变量节点230传递过来的值
wire [5:0] value_check_19_to_variable_230;
wire enable_check_19_to_variable_230;
wire [5:0] value_variable_230_to_check_19;
wire enable_variable_230_to_check_19;
// 对校验节点19的输出值进行拆分
assign value_check_19_to_variable_230 = value_check_19_to_variable[35:30];
assign enable_check_19_to_variable_230 = enable_check_19_to_variable[5];
// 对变量节点230传递过来的值进行组合
assign value_variable_to_check_19[35:30] = value_variable_230_to_check_19;
assign enable_variable_to_check_19[5] = enable_variable_230_to_check_19;


// 校验节点20的接口
wire [35:0] value_variable_to_check_20;
wire [35:0] value_check_20_to_variable;
wire [5:0] enable_variable_to_check_20;
wire [5:0] enable_check_20_to_variable;

// 拆分后校验节点20传递给变量节点17的值以及对变量节点17传递过来的值
wire [5:0] value_check_20_to_variable_17;
wire enable_check_20_to_variable_17;
wire [5:0] value_variable_17_to_check_20;
wire enable_variable_17_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_17 = value_check_20_to_variable[5:0];
assign enable_check_20_to_variable_17 = enable_check_20_to_variable[0];
// 对变量节点17传递过来的值进行组合
assign value_variable_to_check_20[5:0] = value_variable_17_to_check_20;
assign enable_variable_to_check_20[0] = enable_variable_17_to_check_20;

// 拆分后校验节点20传递给变量节点46的值以及对变量节点46传递过来的值
wire [5:0] value_check_20_to_variable_46;
wire enable_check_20_to_variable_46;
wire [5:0] value_variable_46_to_check_20;
wire enable_variable_46_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_46 = value_check_20_to_variable[11:6];
assign enable_check_20_to_variable_46 = enable_check_20_to_variable[1];
// 对变量节点46传递过来的值进行组合
assign value_variable_to_check_20[11:6] = value_variable_46_to_check_20;
assign enable_variable_to_check_20[1] = enable_variable_46_to_check_20;

// 拆分后校验节点20传递给变量节点103的值以及对变量节点103传递过来的值
wire [5:0] value_check_20_to_variable_103;
wire enable_check_20_to_variable_103;
wire [5:0] value_variable_103_to_check_20;
wire enable_variable_103_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_103 = value_check_20_to_variable[17:12];
assign enable_check_20_to_variable_103 = enable_check_20_to_variable[2];
// 对变量节点103传递过来的值进行组合
assign value_variable_to_check_20[17:12] = value_variable_103_to_check_20;
assign enable_variable_to_check_20[2] = enable_variable_103_to_check_20;

// 拆分后校验节点20传递给变量节点147的值以及对变量节点147传递过来的值
wire [5:0] value_check_20_to_variable_147;
wire enable_check_20_to_variable_147;
wire [5:0] value_variable_147_to_check_20;
wire enable_variable_147_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_147 = value_check_20_to_variable[23:18];
assign enable_check_20_to_variable_147 = enable_check_20_to_variable[3];
// 对变量节点147传递过来的值进行组合
assign value_variable_to_check_20[23:18] = value_variable_147_to_check_20;
assign enable_variable_to_check_20[3] = enable_variable_147_to_check_20;

// 拆分后校验节点20传递给变量节点165的值以及对变量节点165传递过来的值
wire [5:0] value_check_20_to_variable_165;
wire enable_check_20_to_variable_165;
wire [5:0] value_variable_165_to_check_20;
wire enable_variable_165_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_165 = value_check_20_to_variable[29:24];
assign enable_check_20_to_variable_165 = enable_check_20_to_variable[4];
// 对变量节点165传递过来的值进行组合
assign value_variable_to_check_20[29:24] = value_variable_165_to_check_20;
assign enable_variable_to_check_20[4] = enable_variable_165_to_check_20;

// 拆分后校验节点20传递给变量节点231的值以及对变量节点231传递过来的值
wire [5:0] value_check_20_to_variable_231;
wire enable_check_20_to_variable_231;
wire [5:0] value_variable_231_to_check_20;
wire enable_variable_231_to_check_20;
// 对校验节点20的输出值进行拆分
assign value_check_20_to_variable_231 = value_check_20_to_variable[35:30];
assign enable_check_20_to_variable_231 = enable_check_20_to_variable[5];
// 对变量节点231传递过来的值进行组合
assign value_variable_to_check_20[35:30] = value_variable_231_to_check_20;
assign enable_variable_to_check_20[5] = enable_variable_231_to_check_20;


// 校验节点21的接口
wire [35:0] value_variable_to_check_21;
wire [35:0] value_check_21_to_variable;
wire [5:0] enable_variable_to_check_21;
wire [5:0] enable_check_21_to_variable;

// 拆分后校验节点21传递给变量节点18的值以及对变量节点18传递过来的值
wire [5:0] value_check_21_to_variable_18;
wire enable_check_21_to_variable_18;
wire [5:0] value_variable_18_to_check_21;
wire enable_variable_18_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_18 = value_check_21_to_variable[5:0];
assign enable_check_21_to_variable_18 = enable_check_21_to_variable[0];
// 对变量节点18传递过来的值进行组合
assign value_variable_to_check_21[5:0] = value_variable_18_to_check_21;
assign enable_variable_to_check_21[0] = enable_variable_18_to_check_21;

// 拆分后校验节点21传递给变量节点61的值以及对变量节点61传递过来的值
wire [5:0] value_check_21_to_variable_61;
wire enable_check_21_to_variable_61;
wire [5:0] value_variable_61_to_check_21;
wire enable_variable_61_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_61 = value_check_21_to_variable[11:6];
assign enable_check_21_to_variable_61 = enable_check_21_to_variable[1];
// 对变量节点61传递过来的值进行组合
assign value_variable_to_check_21[11:6] = value_variable_61_to_check_21;
assign enable_variable_to_check_21[1] = enable_variable_61_to_check_21;

// 拆分后校验节点21传递给变量节点104的值以及对变量节点104传递过来的值
wire [5:0] value_check_21_to_variable_104;
wire enable_check_21_to_variable_104;
wire [5:0] value_variable_104_to_check_21;
wire enable_variable_104_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_104 = value_check_21_to_variable[17:12];
assign enable_check_21_to_variable_104 = enable_check_21_to_variable[2];
// 对变量节点104传递过来的值进行组合
assign value_variable_to_check_21[17:12] = value_variable_104_to_check_21;
assign enable_variable_to_check_21[2] = enable_variable_104_to_check_21;

// 拆分后校验节点21传递给变量节点132的值以及对变量节点132传递过来的值
wire [5:0] value_check_21_to_variable_132;
wire enable_check_21_to_variable_132;
wire [5:0] value_variable_132_to_check_21;
wire enable_variable_132_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_132 = value_check_21_to_variable[23:18];
assign enable_check_21_to_variable_132 = enable_check_21_to_variable[3];
// 对变量节点132传递过来的值进行组合
assign value_variable_to_check_21[23:18] = value_variable_132_to_check_21;
assign enable_variable_to_check_21[3] = enable_variable_132_to_check_21;

// 拆分后校验节点21传递给变量节点188的值以及对变量节点188传递过来的值
wire [5:0] value_check_21_to_variable_188;
wire enable_check_21_to_variable_188;
wire [5:0] value_variable_188_to_check_21;
wire enable_variable_188_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_188 = value_check_21_to_variable[29:24];
assign enable_check_21_to_variable_188 = enable_check_21_to_variable[4];
// 对变量节点188传递过来的值进行组合
assign value_variable_to_check_21[29:24] = value_variable_188_to_check_21;
assign enable_variable_to_check_21[4] = enable_variable_188_to_check_21;

// 拆分后校验节点21传递给变量节点218的值以及对变量节点218传递过来的值
wire [5:0] value_check_21_to_variable_218;
wire enable_check_21_to_variable_218;
wire [5:0] value_variable_218_to_check_21;
wire enable_variable_218_to_check_21;
// 对校验节点21的输出值进行拆分
assign value_check_21_to_variable_218 = value_check_21_to_variable[35:30];
assign enable_check_21_to_variable_218 = enable_check_21_to_variable[5];
// 对变量节点218传递过来的值进行组合
assign value_variable_to_check_21[35:30] = value_variable_218_to_check_21;
assign enable_variable_to_check_21[5] = enable_variable_218_to_check_21;


// 校验节点22的接口
wire [35:0] value_variable_to_check_22;
wire [35:0] value_check_22_to_variable;
wire [5:0] enable_variable_to_check_22;
wire [5:0] enable_check_22_to_variable;

// 拆分后校验节点22传递给变量节点18的值以及对变量节点18传递过来的值
wire [5:0] value_check_22_to_variable_18;
wire enable_check_22_to_variable_18;
wire [5:0] value_variable_18_to_check_22;
wire enable_variable_18_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_18 = value_check_22_to_variable[5:0];
assign enable_check_22_to_variable_18 = enable_check_22_to_variable[0];
// 对变量节点18传递过来的值进行组合
assign value_variable_to_check_22[5:0] = value_variable_18_to_check_22;
assign enable_variable_to_check_22[0] = enable_variable_18_to_check_22;

// 拆分后校验节点22传递给变量节点62的值以及对变量节点62传递过来的值
wire [5:0] value_check_22_to_variable_62;
wire enable_check_22_to_variable_62;
wire [5:0] value_variable_62_to_check_22;
wire enable_variable_62_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_62 = value_check_22_to_variable[11:6];
assign enable_check_22_to_variable_62 = enable_check_22_to_variable[1];
// 对变量节点62传递过来的值进行组合
assign value_variable_to_check_22[11:6] = value_variable_62_to_check_22;
assign enable_variable_to_check_22[1] = enable_variable_62_to_check_22;

// 拆分后校验节点22传递给变量节点96的值以及对变量节点96传递过来的值
wire [5:0] value_check_22_to_variable_96;
wire enable_check_22_to_variable_96;
wire [5:0] value_variable_96_to_check_22;
wire enable_variable_96_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_96 = value_check_22_to_variable[17:12];
assign enable_check_22_to_variable_96 = enable_check_22_to_variable[2];
// 对变量节点96传递过来的值进行组合
assign value_variable_to_check_22[17:12] = value_variable_96_to_check_22;
assign enable_variable_to_check_22[2] = enable_variable_96_to_check_22;

// 拆分后校验节点22传递给变量节点148的值以及对变量节点148传递过来的值
wire [5:0] value_check_22_to_variable_148;
wire enable_check_22_to_variable_148;
wire [5:0] value_variable_148_to_check_22;
wire enable_variable_148_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_148 = value_check_22_to_variable[23:18];
assign enable_check_22_to_variable_148 = enable_check_22_to_variable[3];
// 对变量节点148传递过来的值进行组合
assign value_variable_to_check_22[23:18] = value_variable_148_to_check_22;
assign enable_variable_to_check_22[3] = enable_variable_148_to_check_22;

// 拆分后校验节点22传递给变量节点189的值以及对变量节点189传递过来的值
wire [5:0] value_check_22_to_variable_189;
wire enable_check_22_to_variable_189;
wire [5:0] value_variable_189_to_check_22;
wire enable_variable_189_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_189 = value_check_22_to_variable[29:24];
assign enable_check_22_to_variable_189 = enable_check_22_to_variable[4];
// 对变量节点189传递过来的值进行组合
assign value_variable_to_check_22[29:24] = value_variable_189_to_check_22;
assign enable_variable_to_check_22[4] = enable_variable_189_to_check_22;

// 拆分后校验节点22传递给变量节点226的值以及对变量节点226传递过来的值
wire [5:0] value_check_22_to_variable_226;
wire enable_check_22_to_variable_226;
wire [5:0] value_variable_226_to_check_22;
wire enable_variable_226_to_check_22;
// 对校验节点22的输出值进行拆分
assign value_check_22_to_variable_226 = value_check_22_to_variable[35:30];
assign enable_check_22_to_variable_226 = enable_check_22_to_variable[5];
// 对变量节点226传递过来的值进行组合
assign value_variable_to_check_22[35:30] = value_variable_226_to_check_22;
assign enable_variable_to_check_22[5] = enable_variable_226_to_check_22;


// 校验节点23的接口
wire [35:0] value_variable_to_check_23;
wire [35:0] value_check_23_to_variable;
wire [5:0] enable_variable_to_check_23;
wire [5:0] enable_check_23_to_variable;

// 拆分后校验节点23传递给变量节点19的值以及对变量节点19传递过来的值
wire [5:0] value_check_23_to_variable_19;
wire enable_check_23_to_variable_19;
wire [5:0] value_variable_19_to_check_23;
wire enable_variable_19_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_19 = value_check_23_to_variable[5:0];
assign enable_check_23_to_variable_19 = enable_check_23_to_variable[0];
// 对变量节点19传递过来的值进行组合
assign value_variable_to_check_23[5:0] = value_variable_19_to_check_23;
assign enable_variable_to_check_23[0] = enable_variable_19_to_check_23;

// 拆分后校验节点23传递给变量节点55的值以及对变量节点55传递过来的值
wire [5:0] value_check_23_to_variable_55;
wire enable_check_23_to_variable_55;
wire [5:0] value_variable_55_to_check_23;
wire enable_variable_55_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_55 = value_check_23_to_variable[11:6];
assign enable_check_23_to_variable_55 = enable_check_23_to_variable[1];
// 对变量节点55传递过来的值进行组合
assign value_variable_to_check_23[11:6] = value_variable_55_to_check_23;
assign enable_variable_to_check_23[1] = enable_variable_55_to_check_23;

// 拆分后校验节点23传递给变量节点94的值以及对变量节点94传递过来的值
wire [5:0] value_check_23_to_variable_94;
wire enable_check_23_to_variable_94;
wire [5:0] value_variable_94_to_check_23;
wire enable_variable_94_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_94 = value_check_23_to_variable[17:12];
assign enable_check_23_to_variable_94 = enable_check_23_to_variable[2];
// 对变量节点94传递过来的值进行组合
assign value_variable_to_check_23[17:12] = value_variable_94_to_check_23;
assign enable_variable_to_check_23[2] = enable_variable_94_to_check_23;

// 拆分后校验节点23传递给变量节点149的值以及对变量节点149传递过来的值
wire [5:0] value_check_23_to_variable_149;
wire enable_check_23_to_variable_149;
wire [5:0] value_variable_149_to_check_23;
wire enable_variable_149_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_149 = value_check_23_to_variable[23:18];
assign enable_check_23_to_variable_149 = enable_check_23_to_variable[3];
// 对变量节点149传递过来的值进行组合
assign value_variable_to_check_23[23:18] = value_variable_149_to_check_23;
assign enable_variable_to_check_23[3] = enable_variable_149_to_check_23;

// 拆分后校验节点23传递给变量节点190的值以及对变量节点190传递过来的值
wire [5:0] value_check_23_to_variable_190;
wire enable_check_23_to_variable_190;
wire [5:0] value_variable_190_to_check_23;
wire enable_variable_190_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_190 = value_check_23_to_variable[29:24];
assign enable_check_23_to_variable_190 = enable_check_23_to_variable[4];
// 对变量节点190传递过来的值进行组合
assign value_variable_to_check_23[29:24] = value_variable_190_to_check_23;
assign enable_variable_to_check_23[4] = enable_variable_190_to_check_23;

// 拆分后校验节点23传递给变量节点232的值以及对变量节点232传递过来的值
wire [5:0] value_check_23_to_variable_232;
wire enable_check_23_to_variable_232;
wire [5:0] value_variable_232_to_check_23;
wire enable_variable_232_to_check_23;
// 对校验节点23的输出值进行拆分
assign value_check_23_to_variable_232 = value_check_23_to_variable[35:30];
assign enable_check_23_to_variable_232 = enable_check_23_to_variable[5];
// 对变量节点232传递过来的值进行组合
assign value_variable_to_check_23[35:30] = value_variable_232_to_check_23;
assign enable_variable_to_check_23[5] = enable_variable_232_to_check_23;


// 校验节点24的接口
wire [35:0] value_variable_to_check_24;
wire [35:0] value_check_24_to_variable;
wire [5:0] enable_variable_to_check_24;
wire [5:0] enable_check_24_to_variable;

// 拆分后校验节点24传递给变量节点20的值以及对变量节点20传递过来的值
wire [5:0] value_check_24_to_variable_20;
wire enable_check_24_to_variable_20;
wire [5:0] value_variable_20_to_check_24;
wire enable_variable_20_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_20 = value_check_24_to_variable[5:0];
assign enable_check_24_to_variable_20 = enable_check_24_to_variable[0];
// 对变量节点20传递过来的值进行组合
assign value_variable_to_check_24[5:0] = value_variable_20_to_check_24;
assign enable_variable_to_check_24[0] = enable_variable_20_to_check_24;

// 拆分后校验节点24传递给变量节点61的值以及对变量节点61传递过来的值
wire [5:0] value_check_24_to_variable_61;
wire enable_check_24_to_variable_61;
wire [5:0] value_variable_61_to_check_24;
wire enable_variable_61_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_61 = value_check_24_to_variable[11:6];
assign enable_check_24_to_variable_61 = enable_check_24_to_variable[1];
// 对变量节点61传递过来的值进行组合
assign value_variable_to_check_24[11:6] = value_variable_61_to_check_24;
assign enable_variable_to_check_24[1] = enable_variable_61_to_check_24;

// 拆分后校验节点24传递给变量节点105的值以及对变量节点105传递过来的值
wire [5:0] value_check_24_to_variable_105;
wire enable_check_24_to_variable_105;
wire [5:0] value_variable_105_to_check_24;
wire enable_variable_105_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_105 = value_check_24_to_variable[17:12];
assign enable_check_24_to_variable_105 = enable_check_24_to_variable[2];
// 对变量节点105传递过来的值进行组合
assign value_variable_to_check_24[17:12] = value_variable_105_to_check_24;
assign enable_variable_to_check_24[2] = enable_variable_105_to_check_24;

// 拆分后校验节点24传递给变量节点150的值以及对变量节点150传递过来的值
wire [5:0] value_check_24_to_variable_150;
wire enable_check_24_to_variable_150;
wire [5:0] value_variable_150_to_check_24;
wire enable_variable_150_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_150 = value_check_24_to_variable[23:18];
assign enable_check_24_to_variable_150 = enable_check_24_to_variable[3];
// 对变量节点150传递过来的值进行组合
assign value_variable_to_check_24[23:18] = value_variable_150_to_check_24;
assign enable_variable_to_check_24[3] = enable_variable_150_to_check_24;

// 拆分后校验节点24传递给变量节点182的值以及对变量节点182传递过来的值
wire [5:0] value_check_24_to_variable_182;
wire enable_check_24_to_variable_182;
wire [5:0] value_variable_182_to_check_24;
wire enable_variable_182_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_182 = value_check_24_to_variable[29:24];
assign enable_check_24_to_variable_182 = enable_check_24_to_variable[4];
// 对变量节点182传递过来的值进行组合
assign value_variable_to_check_24[29:24] = value_variable_182_to_check_24;
assign enable_variable_to_check_24[4] = enable_variable_182_to_check_24;

// 拆分后校验节点24传递给变量节点233的值以及对变量节点233传递过来的值
wire [5:0] value_check_24_to_variable_233;
wire enable_check_24_to_variable_233;
wire [5:0] value_variable_233_to_check_24;
wire enable_variable_233_to_check_24;
// 对校验节点24的输出值进行拆分
assign value_check_24_to_variable_233 = value_check_24_to_variable[35:30];
assign enable_check_24_to_variable_233 = enable_check_24_to_variable[5];
// 对变量节点233传递过来的值进行组合
assign value_variable_to_check_24[35:30] = value_variable_233_to_check_24;
assign enable_variable_to_check_24[5] = enable_variable_233_to_check_24;


// 校验节点25的接口
wire [35:0] value_variable_to_check_25;
wire [35:0] value_check_25_to_variable;
wire [5:0] enable_variable_to_check_25;
wire [5:0] enable_check_25_to_variable;

// 拆分后校验节点25传递给变量节点21的值以及对变量节点21传递过来的值
wire [5:0] value_check_25_to_variable_21;
wire enable_check_25_to_variable_21;
wire [5:0] value_variable_21_to_check_25;
wire enable_variable_21_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_21 = value_check_25_to_variable[5:0];
assign enable_check_25_to_variable_21 = enable_check_25_to_variable[0];
// 对变量节点21传递过来的值进行组合
assign value_variable_to_check_25[5:0] = value_variable_21_to_check_25;
assign enable_variable_to_check_25[0] = enable_variable_21_to_check_25;

// 拆分后校验节点25传递给变量节点50的值以及对变量节点50传递过来的值
wire [5:0] value_check_25_to_variable_50;
wire enable_check_25_to_variable_50;
wire [5:0] value_variable_50_to_check_25;
wire enable_variable_50_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_50 = value_check_25_to_variable[11:6];
assign enable_check_25_to_variable_50 = enable_check_25_to_variable[1];
// 对变量节点50传递过来的值进行组合
assign value_variable_to_check_25[11:6] = value_variable_50_to_check_25;
assign enable_variable_to_check_25[1] = enable_variable_50_to_check_25;

// 拆分后校验节点25传递给变量节点106的值以及对变量节点106传递过来的值
wire [5:0] value_check_25_to_variable_106;
wire enable_check_25_to_variable_106;
wire [5:0] value_variable_106_to_check_25;
wire enable_variable_106_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_106 = value_check_25_to_variable[17:12];
assign enable_check_25_to_variable_106 = enable_check_25_to_variable[2];
// 对变量节点106传递过来的值进行组合
assign value_variable_to_check_25[17:12] = value_variable_106_to_check_25;
assign enable_variable_to_check_25[2] = enable_variable_106_to_check_25;

// 拆分后校验节点25传递给变量节点137的值以及对变量节点137传递过来的值
wire [5:0] value_check_25_to_variable_137;
wire enable_check_25_to_variable_137;
wire [5:0] value_variable_137_to_check_25;
wire enable_variable_137_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_137 = value_check_25_to_variable[23:18];
assign enable_check_25_to_variable_137 = enable_check_25_to_variable[3];
// 对变量节点137传递过来的值进行组合
assign value_variable_to_check_25[23:18] = value_variable_137_to_check_25;
assign enable_variable_to_check_25[3] = enable_variable_137_to_check_25;

// 拆分后校验节点25传递给变量节点191的值以及对变量节点191传递过来的值
wire [5:0] value_check_25_to_variable_191;
wire enable_check_25_to_variable_191;
wire [5:0] value_variable_191_to_check_25;
wire enable_variable_191_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_191 = value_check_25_to_variable[29:24];
assign enable_check_25_to_variable_191 = enable_check_25_to_variable[4];
// 对变量节点191传递过来的值进行组合
assign value_variable_to_check_25[29:24] = value_variable_191_to_check_25;
assign enable_variable_to_check_25[4] = enable_variable_191_to_check_25;

// 拆分后校验节点25传递给变量节点234的值以及对变量节点234传递过来的值
wire [5:0] value_check_25_to_variable_234;
wire enable_check_25_to_variable_234;
wire [5:0] value_variable_234_to_check_25;
wire enable_variable_234_to_check_25;
// 对校验节点25的输出值进行拆分
assign value_check_25_to_variable_234 = value_check_25_to_variable[35:30];
assign enable_check_25_to_variable_234 = enable_check_25_to_variable[5];
// 对变量节点234传递过来的值进行组合
assign value_variable_to_check_25[35:30] = value_variable_234_to_check_25;
assign enable_variable_to_check_25[5] = enable_variable_234_to_check_25;


// 校验节点26的接口
wire [35:0] value_variable_to_check_26;
wire [35:0] value_check_26_to_variable;
wire [5:0] enable_variable_to_check_26;
wire [5:0] enable_check_26_to_variable;

// 拆分后校验节点26传递给变量节点22的值以及对变量节点22传递过来的值
wire [5:0] value_check_26_to_variable_22;
wire enable_check_26_to_variable_22;
wire [5:0] value_variable_22_to_check_26;
wire enable_variable_22_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_22 = value_check_26_to_variable[5:0];
assign enable_check_26_to_variable_22 = enable_check_26_to_variable[0];
// 对变量节点22传递过来的值进行组合
assign value_variable_to_check_26[5:0] = value_variable_22_to_check_26;
assign enable_variable_to_check_26[0] = enable_variable_22_to_check_26;

// 拆分后校验节点26传递给变量节点63的值以及对变量节点63传递过来的值
wire [5:0] value_check_26_to_variable_63;
wire enable_check_26_to_variable_63;
wire [5:0] value_variable_63_to_check_26;
wire enable_variable_63_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_63 = value_check_26_to_variable[11:6];
assign enable_check_26_to_variable_63 = enable_check_26_to_variable[1];
// 对变量节点63传递过来的值进行组合
assign value_variable_to_check_26[11:6] = value_variable_63_to_check_26;
assign enable_variable_to_check_26[1] = enable_variable_63_to_check_26;

// 拆分后校验节点26传递给变量节点95的值以及对变量节点95传递过来的值
wire [5:0] value_check_26_to_variable_95;
wire enable_check_26_to_variable_95;
wire [5:0] value_variable_95_to_check_26;
wire enable_variable_95_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_95 = value_check_26_to_variable[17:12];
assign enable_check_26_to_variable_95 = enable_check_26_to_variable[2];
// 对变量节点95传递过来的值进行组合
assign value_variable_to_check_26[17:12] = value_variable_95_to_check_26;
assign enable_variable_to_check_26[2] = enable_variable_95_to_check_26;

// 拆分后校验节点26传递给变量节点151的值以及对变量节点151传递过来的值
wire [5:0] value_check_26_to_variable_151;
wire enable_check_26_to_variable_151;
wire [5:0] value_variable_151_to_check_26;
wire enable_variable_151_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_151 = value_check_26_to_variable[23:18];
assign enable_check_26_to_variable_151 = enable_check_26_to_variable[3];
// 对变量节点151传递过来的值进行组合
assign value_variable_to_check_26[23:18] = value_variable_151_to_check_26;
assign enable_variable_to_check_26[3] = enable_variable_151_to_check_26;

// 拆分后校验节点26传递给变量节点192的值以及对变量节点192传递过来的值
wire [5:0] value_check_26_to_variable_192;
wire enable_check_26_to_variable_192;
wire [5:0] value_variable_192_to_check_26;
wire enable_variable_192_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_192 = value_check_26_to_variable[29:24];
assign enable_check_26_to_variable_192 = enable_check_26_to_variable[4];
// 对变量节点192传递过来的值进行组合
assign value_variable_to_check_26[29:24] = value_variable_192_to_check_26;
assign enable_variable_to_check_26[4] = enable_variable_192_to_check_26;

// 拆分后校验节点26传递给变量节点235的值以及对变量节点235传递过来的值
wire [5:0] value_check_26_to_variable_235;
wire enable_check_26_to_variable_235;
wire [5:0] value_variable_235_to_check_26;
wire enable_variable_235_to_check_26;
// 对校验节点26的输出值进行拆分
assign value_check_26_to_variable_235 = value_check_26_to_variable[35:30];
assign enable_check_26_to_variable_235 = enable_check_26_to_variable[5];
// 对变量节点235传递过来的值进行组合
assign value_variable_to_check_26[35:30] = value_variable_235_to_check_26;
assign enable_variable_to_check_26[5] = enable_variable_235_to_check_26;


// 校验节点27的接口
wire [35:0] value_variable_to_check_27;
wire [35:0] value_check_27_to_variable;
wire [5:0] enable_variable_to_check_27;
wire [5:0] enable_check_27_to_variable;

// 拆分后校验节点27传递给变量节点23的值以及对变量节点23传递过来的值
wire [5:0] value_check_27_to_variable_23;
wire enable_check_27_to_variable_23;
wire [5:0] value_variable_23_to_check_27;
wire enable_variable_23_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_23 = value_check_27_to_variable[5:0];
assign enable_check_27_to_variable_23 = enable_check_27_to_variable[0];
// 对变量节点23传递过来的值进行组合
assign value_variable_to_check_27[5:0] = value_variable_23_to_check_27;
assign enable_variable_to_check_27[0] = enable_variable_23_to_check_27;

// 拆分后校验节点27传递给变量节点64的值以及对变量节点64传递过来的值
wire [5:0] value_check_27_to_variable_64;
wire enable_check_27_to_variable_64;
wire [5:0] value_variable_64_to_check_27;
wire enable_variable_64_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_64 = value_check_27_to_variable[11:6];
assign enable_check_27_to_variable_64 = enable_check_27_to_variable[1];
// 对变量节点64传递过来的值进行组合
assign value_variable_to_check_27[11:6] = value_variable_64_to_check_27;
assign enable_variable_to_check_27[1] = enable_variable_64_to_check_27;

// 拆分后校验节点27传递给变量节点107的值以及对变量节点107传递过来的值
wire [5:0] value_check_27_to_variable_107;
wire enable_check_27_to_variable_107;
wire [5:0] value_variable_107_to_check_27;
wire enable_variable_107_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_107 = value_check_27_to_variable[17:12];
assign enable_check_27_to_variable_107 = enable_check_27_to_variable[2];
// 对变量节点107传递过来的值进行组合
assign value_variable_to_check_27[17:12] = value_variable_107_to_check_27;
assign enable_variable_to_check_27[2] = enable_variable_107_to_check_27;

// 拆分后校验节点27传递给变量节点152的值以及对变量节点152传递过来的值
wire [5:0] value_check_27_to_variable_152;
wire enable_check_27_to_variable_152;
wire [5:0] value_variable_152_to_check_27;
wire enable_variable_152_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_152 = value_check_27_to_variable[23:18];
assign enable_check_27_to_variable_152 = enable_check_27_to_variable[3];
// 对变量节点152传递过来的值进行组合
assign value_variable_to_check_27[23:18] = value_variable_152_to_check_27;
assign enable_variable_to_check_27[3] = enable_variable_152_to_check_27;

// 拆分后校验节点27传递给变量节点193的值以及对变量节点193传递过来的值
wire [5:0] value_check_27_to_variable_193;
wire enable_check_27_to_variable_193;
wire [5:0] value_variable_193_to_check_27;
wire enable_variable_193_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_193 = value_check_27_to_variable[29:24];
assign enable_check_27_to_variable_193 = enable_check_27_to_variable[4];
// 对变量节点193传递过来的值进行组合
assign value_variable_to_check_27[29:24] = value_variable_193_to_check_27;
assign enable_variable_to_check_27[4] = enable_variable_193_to_check_27;

// 拆分后校验节点27传递给变量节点225的值以及对变量节点225传递过来的值
wire [5:0] value_check_27_to_variable_225;
wire enable_check_27_to_variable_225;
wire [5:0] value_variable_225_to_check_27;
wire enable_variable_225_to_check_27;
// 对校验节点27的输出值进行拆分
assign value_check_27_to_variable_225 = value_check_27_to_variable[35:30];
assign enable_check_27_to_variable_225 = enable_check_27_to_variable[5];
// 对变量节点225传递过来的值进行组合
assign value_variable_to_check_27[35:30] = value_variable_225_to_check_27;
assign enable_variable_to_check_27[5] = enable_variable_225_to_check_27;


// 校验节点28的接口
wire [35:0] value_variable_to_check_28;
wire [35:0] value_check_28_to_variable;
wire [5:0] enable_variable_to_check_28;
wire [5:0] enable_check_28_to_variable;

// 拆分后校验节点28传递给变量节点24的值以及对变量节点24传递过来的值
wire [5:0] value_check_28_to_variable_24;
wire enable_check_28_to_variable_24;
wire [5:0] value_variable_24_to_check_28;
wire enable_variable_24_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_24 = value_check_28_to_variable[5:0];
assign enable_check_28_to_variable_24 = enable_check_28_to_variable[0];
// 对变量节点24传递过来的值进行组合
assign value_variable_to_check_28[5:0] = value_variable_24_to_check_28;
assign enable_variable_to_check_28[0] = enable_variable_24_to_check_28;

// 拆分后校验节点28传递给变量节点65的值以及对变量节点65传递过来的值
wire [5:0] value_check_28_to_variable_65;
wire enable_check_28_to_variable_65;
wire [5:0] value_variable_65_to_check_28;
wire enable_variable_65_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_65 = value_check_28_to_variable[11:6];
assign enable_check_28_to_variable_65 = enable_check_28_to_variable[1];
// 对变量节点65传递过来的值进行组合
assign value_variable_to_check_28[11:6] = value_variable_65_to_check_28;
assign enable_variable_to_check_28[1] = enable_variable_65_to_check_28;

// 拆分后校验节点28传递给变量节点89的值以及对变量节点89传递过来的值
wire [5:0] value_check_28_to_variable_89;
wire enable_check_28_to_variable_89;
wire [5:0] value_variable_89_to_check_28;
wire enable_variable_89_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_89 = value_check_28_to_variable[17:12];
assign enable_check_28_to_variable_89 = enable_check_28_to_variable[2];
// 对变量节点89传递过来的值进行组合
assign value_variable_to_check_28[17:12] = value_variable_89_to_check_28;
assign enable_variable_to_check_28[2] = enable_variable_89_to_check_28;

// 拆分后校验节点28传递给变量节点153的值以及对变量节点153传递过来的值
wire [5:0] value_check_28_to_variable_153;
wire enable_check_28_to_variable_153;
wire [5:0] value_variable_153_to_check_28;
wire enable_variable_153_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_153 = value_check_28_to_variable[23:18];
assign enable_check_28_to_variable_153 = enable_check_28_to_variable[3];
// 对变量节点153传递过来的值进行组合
assign value_variable_to_check_28[23:18] = value_variable_153_to_check_28;
assign enable_variable_to_check_28[3] = enable_variable_153_to_check_28;

// 拆分后校验节点28传递给变量节点194的值以及对变量节点194传递过来的值
wire [5:0] value_check_28_to_variable_194;
wire enable_check_28_to_variable_194;
wire [5:0] value_variable_194_to_check_28;
wire enable_variable_194_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_194 = value_check_28_to_variable[29:24];
assign enable_check_28_to_variable_194 = enable_check_28_to_variable[4];
// 对变量节点194传递过来的值进行组合
assign value_variable_to_check_28[29:24] = value_variable_194_to_check_28;
assign enable_variable_to_check_28[4] = enable_variable_194_to_check_28;

// 拆分后校验节点28传递给变量节点236的值以及对变量节点236传递过来的值
wire [5:0] value_check_28_to_variable_236;
wire enable_check_28_to_variable_236;
wire [5:0] value_variable_236_to_check_28;
wire enable_variable_236_to_check_28;
// 对校验节点28的输出值进行拆分
assign value_check_28_to_variable_236 = value_check_28_to_variable[35:30];
assign enable_check_28_to_variable_236 = enable_check_28_to_variable[5];
// 对变量节点236传递过来的值进行组合
assign value_variable_to_check_28[35:30] = value_variable_236_to_check_28;
assign enable_variable_to_check_28[5] = enable_variable_236_to_check_28;


// 校验节点29的接口
wire [35:0] value_variable_to_check_29;
wire [35:0] value_check_29_to_variable;
wire [5:0] enable_variable_to_check_29;
wire [5:0] enable_check_29_to_variable;

// 拆分后校验节点29传递给变量节点11的值以及对变量节点11传递过来的值
wire [5:0] value_check_29_to_variable_11;
wire enable_check_29_to_variable_11;
wire [5:0] value_variable_11_to_check_29;
wire enable_variable_11_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_11 = value_check_29_to_variable[5:0];
assign enable_check_29_to_variable_11 = enable_check_29_to_variable[0];
// 对变量节点11传递过来的值进行组合
assign value_variable_to_check_29[5:0] = value_variable_11_to_check_29;
assign enable_variable_to_check_29[0] = enable_variable_11_to_check_29;

// 拆分后校验节点29传递给变量节点66的值以及对变量节点66传递过来的值
wire [5:0] value_check_29_to_variable_66;
wire enable_check_29_to_variable_66;
wire [5:0] value_variable_66_to_check_29;
wire enable_variable_66_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_66 = value_check_29_to_variable[11:6];
assign enable_check_29_to_variable_66 = enable_check_29_to_variable[1];
// 对变量节点66传递过来的值进行组合
assign value_variable_to_check_29[11:6] = value_variable_66_to_check_29;
assign enable_variable_to_check_29[1] = enable_variable_66_to_check_29;

// 拆分后校验节点29传递给变量节点104的值以及对变量节点104传递过来的值
wire [5:0] value_check_29_to_variable_104;
wire enable_check_29_to_variable_104;
wire [5:0] value_variable_104_to_check_29;
wire enable_variable_104_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_104 = value_check_29_to_variable[17:12];
assign enable_check_29_to_variable_104 = enable_check_29_to_variable[2];
// 对变量节点104传递过来的值进行组合
assign value_variable_to_check_29[17:12] = value_variable_104_to_check_29;
assign enable_variable_to_check_29[2] = enable_variable_104_to_check_29;

// 拆分后校验节点29传递给变量节点154的值以及对变量节点154传递过来的值
wire [5:0] value_check_29_to_variable_154;
wire enable_check_29_to_variable_154;
wire [5:0] value_variable_154_to_check_29;
wire enable_variable_154_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_154 = value_check_29_to_variable[23:18];
assign enable_check_29_to_variable_154 = enable_check_29_to_variable[3];
// 对变量节点154传递过来的值进行组合
assign value_variable_to_check_29[23:18] = value_variable_154_to_check_29;
assign enable_variable_to_check_29[3] = enable_variable_154_to_check_29;

// 拆分后校验节点29传递给变量节点180的值以及对变量节点180传递过来的值
wire [5:0] value_check_29_to_variable_180;
wire enable_check_29_to_variable_180;
wire [5:0] value_variable_180_to_check_29;
wire enable_variable_180_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_180 = value_check_29_to_variable[29:24];
assign enable_check_29_to_variable_180 = enable_check_29_to_variable[4];
// 对变量节点180传递过来的值进行组合
assign value_variable_to_check_29[29:24] = value_variable_180_to_check_29;
assign enable_variable_to_check_29[4] = enable_variable_180_to_check_29;

// 拆分后校验节点29传递给变量节点237的值以及对变量节点237传递过来的值
wire [5:0] value_check_29_to_variable_237;
wire enable_check_29_to_variable_237;
wire [5:0] value_variable_237_to_check_29;
wire enable_variable_237_to_check_29;
// 对校验节点29的输出值进行拆分
assign value_check_29_to_variable_237 = value_check_29_to_variable[35:30];
assign enable_check_29_to_variable_237 = enable_check_29_to_variable[5];
// 对变量节点237传递过来的值进行组合
assign value_variable_to_check_29[35:30] = value_variable_237_to_check_29;
assign enable_variable_to_check_29[5] = enable_variable_237_to_check_29;


// 校验节点30的接口
wire [35:0] value_variable_to_check_30;
wire [35:0] value_check_30_to_variable;
wire [5:0] enable_variable_to_check_30;
wire [5:0] enable_check_30_to_variable;

// 拆分后校验节点30传递给变量节点25的值以及对变量节点25传递过来的值
wire [5:0] value_check_30_to_variable_25;
wire enable_check_30_to_variable_25;
wire [5:0] value_variable_25_to_check_30;
wire enable_variable_25_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_25 = value_check_30_to_variable[5:0];
assign enable_check_30_to_variable_25 = enable_check_30_to_variable[0];
// 对变量节点25传递过来的值进行组合
assign value_variable_to_check_30[5:0] = value_variable_25_to_check_30;
assign enable_variable_to_check_30[0] = enable_variable_25_to_check_30;

// 拆分后校验节点30传递给变量节点57的值以及对变量节点57传递过来的值
wire [5:0] value_check_30_to_variable_57;
wire enable_check_30_to_variable_57;
wire [5:0] value_variable_57_to_check_30;
wire enable_variable_57_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_57 = value_check_30_to_variable[11:6];
assign enable_check_30_to_variable_57 = enable_check_30_to_variable[1];
// 对变量节点57传递过来的值进行组合
assign value_variable_to_check_30[11:6] = value_variable_57_to_check_30;
assign enable_variable_to_check_30[1] = enable_variable_57_to_check_30;

// 拆分后校验节点30传递给变量节点108的值以及对变量节点108传递过来的值
wire [5:0] value_check_30_to_variable_108;
wire enable_check_30_to_variable_108;
wire [5:0] value_variable_108_to_check_30;
wire enable_variable_108_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_108 = value_check_30_to_variable[17:12];
assign enable_check_30_to_variable_108 = enable_check_30_to_variable[2];
// 对变量节点108传递过来的值进行组合
assign value_variable_to_check_30[17:12] = value_variable_108_to_check_30;
assign enable_variable_to_check_30[2] = enable_variable_108_to_check_30;

// 拆分后校验节点30传递给变量节点155的值以及对变量节点155传递过来的值
wire [5:0] value_check_30_to_variable_155;
wire enable_check_30_to_variable_155;
wire [5:0] value_variable_155_to_check_30;
wire enable_variable_155_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_155 = value_check_30_to_variable[23:18];
assign enable_check_30_to_variable_155 = enable_check_30_to_variable[3];
// 对变量节点155传递过来的值进行组合
assign value_variable_to_check_30[23:18] = value_variable_155_to_check_30;
assign enable_variable_to_check_30[3] = enable_variable_155_to_check_30;

// 拆分后校验节点30传递给变量节点195的值以及对变量节点195传递过来的值
wire [5:0] value_check_30_to_variable_195;
wire enable_check_30_to_variable_195;
wire [5:0] value_variable_195_to_check_30;
wire enable_variable_195_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_195 = value_check_30_to_variable[29:24];
assign enable_check_30_to_variable_195 = enable_check_30_to_variable[4];
// 对变量节点195传递过来的值进行组合
assign value_variable_to_check_30[29:24] = value_variable_195_to_check_30;
assign enable_variable_to_check_30[4] = enable_variable_195_to_check_30;

// 拆分后校验节点30传递给变量节点220的值以及对变量节点220传递过来的值
wire [5:0] value_check_30_to_variable_220;
wire enable_check_30_to_variable_220;
wire [5:0] value_variable_220_to_check_30;
wire enable_variable_220_to_check_30;
// 对校验节点30的输出值进行拆分
assign value_check_30_to_variable_220 = value_check_30_to_variable[35:30];
assign enable_check_30_to_variable_220 = enable_check_30_to_variable[5];
// 对变量节点220传递过来的值进行组合
assign value_variable_to_check_30[35:30] = value_variable_220_to_check_30;
assign enable_variable_to_check_30[5] = enable_variable_220_to_check_30;


// 校验节点31的接口
wire [35:0] value_variable_to_check_31;
wire [35:0] value_check_31_to_variable;
wire [5:0] enable_variable_to_check_31;
wire [5:0] enable_check_31_to_variable;

// 拆分后校验节点31传递给变量节点26的值以及对变量节点26传递过来的值
wire [5:0] value_check_31_to_variable_26;
wire enable_check_31_to_variable_26;
wire [5:0] value_variable_26_to_check_31;
wire enable_variable_26_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_26 = value_check_31_to_variable[5:0];
assign enable_check_31_to_variable_26 = enable_check_31_to_variable[0];
// 对变量节点26传递过来的值进行组合
assign value_variable_to_check_31[5:0] = value_variable_26_to_check_31;
assign enable_variable_to_check_31[0] = enable_variable_26_to_check_31;

// 拆分后校验节点31传递给变量节点59的值以及对变量节点59传递过来的值
wire [5:0] value_check_31_to_variable_59;
wire enable_check_31_to_variable_59;
wire [5:0] value_variable_59_to_check_31;
wire enable_variable_59_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_59 = value_check_31_to_variable[11:6];
assign enable_check_31_to_variable_59 = enable_check_31_to_variable[1];
// 对变量节点59传递过来的值进行组合
assign value_variable_to_check_31[11:6] = value_variable_59_to_check_31;
assign enable_variable_to_check_31[1] = enable_variable_59_to_check_31;

// 拆分后校验节点31传递给变量节点109的值以及对变量节点109传递过来的值
wire [5:0] value_check_31_to_variable_109;
wire enable_check_31_to_variable_109;
wire [5:0] value_variable_109_to_check_31;
wire enable_variable_109_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_109 = value_check_31_to_variable[17:12];
assign enable_check_31_to_variable_109 = enable_check_31_to_variable[2];
// 对变量节点109传递过来的值进行组合
assign value_variable_to_check_31[17:12] = value_variable_109_to_check_31;
assign enable_variable_to_check_31[2] = enable_variable_109_to_check_31;

// 拆分后校验节点31传递给变量节点156的值以及对变量节点156传递过来的值
wire [5:0] value_check_31_to_variable_156;
wire enable_check_31_to_variable_156;
wire [5:0] value_variable_156_to_check_31;
wire enable_variable_156_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_156 = value_check_31_to_variable[23:18];
assign enable_check_31_to_variable_156 = enable_check_31_to_variable[3];
// 对变量节点156传递过来的值进行组合
assign value_variable_to_check_31[23:18] = value_variable_156_to_check_31;
assign enable_variable_to_check_31[3] = enable_variable_156_to_check_31;

// 拆分后校验节点31传递给变量节点195的值以及对变量节点195传递过来的值
wire [5:0] value_check_31_to_variable_195;
wire enable_check_31_to_variable_195;
wire [5:0] value_variable_195_to_check_31;
wire enable_variable_195_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_195 = value_check_31_to_variable[29:24];
assign enable_check_31_to_variable_195 = enable_check_31_to_variable[4];
// 对变量节点195传递过来的值进行组合
assign value_variable_to_check_31[29:24] = value_variable_195_to_check_31;
assign enable_variable_to_check_31[4] = enable_variable_195_to_check_31;

// 拆分后校验节点31传递给变量节点236的值以及对变量节点236传递过来的值
wire [5:0] value_check_31_to_variable_236;
wire enable_check_31_to_variable_236;
wire [5:0] value_variable_236_to_check_31;
wire enable_variable_236_to_check_31;
// 对校验节点31的输出值进行拆分
assign value_check_31_to_variable_236 = value_check_31_to_variable[35:30];
assign enable_check_31_to_variable_236 = enable_check_31_to_variable[5];
// 对变量节点236传递过来的值进行组合
assign value_variable_to_check_31[35:30] = value_variable_236_to_check_31;
assign enable_variable_to_check_31[5] = enable_variable_236_to_check_31;


// 校验节点32的接口
wire [35:0] value_variable_to_check_32;
wire [35:0] value_check_32_to_variable;
wire [5:0] enable_variable_to_check_32;
wire [5:0] enable_check_32_to_variable;

// 拆分后校验节点32传递给变量节点27的值以及对变量节点27传递过来的值
wire [5:0] value_check_32_to_variable_27;
wire enable_check_32_to_variable_27;
wire [5:0] value_variable_27_to_check_32;
wire enable_variable_27_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_27 = value_check_32_to_variable[5:0];
assign enable_check_32_to_variable_27 = enable_check_32_to_variable[0];
// 对变量节点27传递过来的值进行组合
assign value_variable_to_check_32[5:0] = value_variable_27_to_check_32;
assign enable_variable_to_check_32[0] = enable_variable_27_to_check_32;

// 拆分后校验节点32传递给变量节点67的值以及对变量节点67传递过来的值
wire [5:0] value_check_32_to_variable_67;
wire enable_check_32_to_variable_67;
wire [5:0] value_variable_67_to_check_32;
wire enable_variable_67_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_67 = value_check_32_to_variable[11:6];
assign enable_check_32_to_variable_67 = enable_check_32_to_variable[1];
// 对变量节点67传递过来的值进行组合
assign value_variable_to_check_32[11:6] = value_variable_67_to_check_32;
assign enable_variable_to_check_32[1] = enable_variable_67_to_check_32;

// 拆分后校验节点32传递给变量节点110的值以及对变量节点110传递过来的值
wire [5:0] value_check_32_to_variable_110;
wire enable_check_32_to_variable_110;
wire [5:0] value_variable_110_to_check_32;
wire enable_variable_110_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_110 = value_check_32_to_variable[17:12];
assign enable_check_32_to_variable_110 = enable_check_32_to_variable[2];
// 对变量节点110传递过来的值进行组合
assign value_variable_to_check_32[17:12] = value_variable_110_to_check_32;
assign enable_variable_to_check_32[2] = enable_variable_110_to_check_32;

// 拆分后校验节点32传递给变量节点157的值以及对变量节点157传递过来的值
wire [5:0] value_check_32_to_variable_157;
wire enable_check_32_to_variable_157;
wire [5:0] value_variable_157_to_check_32;
wire enable_variable_157_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_157 = value_check_32_to_variable[23:18];
assign enable_check_32_to_variable_157 = enable_check_32_to_variable[3];
// 对变量节点157传递过来的值进行组合
assign value_variable_to_check_32[23:18] = value_variable_157_to_check_32;
assign enable_variable_to_check_32[3] = enable_variable_157_to_check_32;

// 拆分后校验节点32传递给变量节点196的值以及对变量节点196传递过来的值
wire [5:0] value_check_32_to_variable_196;
wire enable_check_32_to_variable_196;
wire [5:0] value_variable_196_to_check_32;
wire enable_variable_196_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_196 = value_check_32_to_variable[29:24];
assign enable_check_32_to_variable_196 = enable_check_32_to_variable[4];
// 对变量节点196传递过来的值进行组合
assign value_variable_to_check_32[29:24] = value_variable_196_to_check_32;
assign enable_variable_to_check_32[4] = enable_variable_196_to_check_32;

// 拆分后校验节点32传递给变量节点214的值以及对变量节点214传递过来的值
wire [5:0] value_check_32_to_variable_214;
wire enable_check_32_to_variable_214;
wire [5:0] value_variable_214_to_check_32;
wire enable_variable_214_to_check_32;
// 对校验节点32的输出值进行拆分
assign value_check_32_to_variable_214 = value_check_32_to_variable[35:30];
assign enable_check_32_to_variable_214 = enable_check_32_to_variable[5];
// 对变量节点214传递过来的值进行组合
assign value_variable_to_check_32[35:30] = value_variable_214_to_check_32;
assign enable_variable_to_check_32[5] = enable_variable_214_to_check_32;


// 校验节点33的接口
wire [35:0] value_variable_to_check_33;
wire [35:0] value_check_33_to_variable;
wire [5:0] enable_variable_to_check_33;
wire [5:0] enable_check_33_to_variable;

// 拆分后校验节点33传递给变量节点28的值以及对变量节点28传递过来的值
wire [5:0] value_check_33_to_variable_28;
wire enable_check_33_to_variable_28;
wire [5:0] value_variable_28_to_check_33;
wire enable_variable_28_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_28 = value_check_33_to_variable[5:0];
assign enable_check_33_to_variable_28 = enable_check_33_to_variable[0];
// 对变量节点28传递过来的值进行组合
assign value_variable_to_check_33[5:0] = value_variable_28_to_check_33;
assign enable_variable_to_check_33[0] = enable_variable_28_to_check_33;

// 拆分后校验节点33传递给变量节点49的值以及对变量节点49传递过来的值
wire [5:0] value_check_33_to_variable_49;
wire enable_check_33_to_variable_49;
wire [5:0] value_variable_49_to_check_33;
wire enable_variable_49_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_49 = value_check_33_to_variable[11:6];
assign enable_check_33_to_variable_49 = enable_check_33_to_variable[1];
// 对变量节点49传递过来的值进行组合
assign value_variable_to_check_33[11:6] = value_variable_49_to_check_33;
assign enable_variable_to_check_33[1] = enable_variable_49_to_check_33;

// 拆分后校验节点33传递给变量节点111的值以及对变量节点111传递过来的值
wire [5:0] value_check_33_to_variable_111;
wire enable_check_33_to_variable_111;
wire [5:0] value_variable_111_to_check_33;
wire enable_variable_111_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_111 = value_check_33_to_variable[17:12];
assign enable_check_33_to_variable_111 = enable_check_33_to_variable[2];
// 对变量节点111传递过来的值进行组合
assign value_variable_to_check_33[17:12] = value_variable_111_to_check_33;
assign enable_variable_to_check_33[2] = enable_variable_111_to_check_33;

// 拆分后校验节点33传递给变量节点158的值以及对变量节点158传递过来的值
wire [5:0] value_check_33_to_variable_158;
wire enable_check_33_to_variable_158;
wire [5:0] value_variable_158_to_check_33;
wire enable_variable_158_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_158 = value_check_33_to_variable[23:18];
assign enable_check_33_to_variable_158 = enable_check_33_to_variable[3];
// 对变量节点158传递过来的值进行组合
assign value_variable_to_check_33[23:18] = value_variable_158_to_check_33;
assign enable_variable_to_check_33[3] = enable_variable_158_to_check_33;

// 拆分后校验节点33传递给变量节点189的值以及对变量节点189传递过来的值
wire [5:0] value_check_33_to_variable_189;
wire enable_check_33_to_variable_189;
wire [5:0] value_variable_189_to_check_33;
wire enable_variable_189_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_189 = value_check_33_to_variable[29:24];
assign enable_check_33_to_variable_189 = enable_check_33_to_variable[4];
// 对变量节点189传递过来的值进行组合
assign value_variable_to_check_33[29:24] = value_variable_189_to_check_33;
assign enable_variable_to_check_33[4] = enable_variable_189_to_check_33;

// 拆分后校验节点33传递给变量节点225的值以及对变量节点225传递过来的值
wire [5:0] value_check_33_to_variable_225;
wire enable_check_33_to_variable_225;
wire [5:0] value_variable_225_to_check_33;
wire enable_variable_225_to_check_33;
// 对校验节点33的输出值进行拆分
assign value_check_33_to_variable_225 = value_check_33_to_variable[35:30];
assign enable_check_33_to_variable_225 = enable_check_33_to_variable[5];
// 对变量节点225传递过来的值进行组合
assign value_variable_to_check_33[35:30] = value_variable_225_to_check_33;
assign enable_variable_to_check_33[5] = enable_variable_225_to_check_33;


// 校验节点34的接口
wire [35:0] value_variable_to_check_34;
wire [35:0] value_check_34_to_variable;
wire [5:0] enable_variable_to_check_34;
wire [5:0] enable_check_34_to_variable;

// 拆分后校验节点34传递给变量节点17的值以及对变量节点17传递过来的值
wire [5:0] value_check_34_to_variable_17;
wire enable_check_34_to_variable_17;
wire [5:0] value_variable_17_to_check_34;
wire enable_variable_17_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_17 = value_check_34_to_variable[5:0];
assign enable_check_34_to_variable_17 = enable_check_34_to_variable[0];
// 对变量节点17传递过来的值进行组合
assign value_variable_to_check_34[5:0] = value_variable_17_to_check_34;
assign enable_variable_to_check_34[0] = enable_variable_17_to_check_34;

// 拆分后校验节点34传递给变量节点52的值以及对变量节点52传递过来的值
wire [5:0] value_check_34_to_variable_52;
wire enable_check_34_to_variable_52;
wire [5:0] value_variable_52_to_check_34;
wire enable_variable_52_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_52 = value_check_34_to_variable[11:6];
assign enable_check_34_to_variable_52 = enable_check_34_to_variable[1];
// 对变量节点52传递过来的值进行组合
assign value_variable_to_check_34[11:6] = value_variable_52_to_check_34;
assign enable_variable_to_check_34[1] = enable_variable_52_to_check_34;

// 拆分后校验节点34传递给变量节点112的值以及对变量节点112传递过来的值
wire [5:0] value_check_34_to_variable_112;
wire enable_check_34_to_variable_112;
wire [5:0] value_variable_112_to_check_34;
wire enable_variable_112_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_112 = value_check_34_to_variable[17:12];
assign enable_check_34_to_variable_112 = enable_check_34_to_variable[2];
// 对变量节点112传递过来的值进行组合
assign value_variable_to_check_34[17:12] = value_variable_112_to_check_34;
assign enable_variable_to_check_34[2] = enable_variable_112_to_check_34;

// 拆分后校验节点34传递给变量节点135的值以及对变量节点135传递过来的值
wire [5:0] value_check_34_to_variable_135;
wire enable_check_34_to_variable_135;
wire [5:0] value_variable_135_to_check_34;
wire enable_variable_135_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_135 = value_check_34_to_variable[23:18];
assign enable_check_34_to_variable_135 = enable_check_34_to_variable[3];
// 对变量节点135传递过来的值进行组合
assign value_variable_to_check_34[23:18] = value_variable_135_to_check_34;
assign enable_variable_to_check_34[3] = enable_variable_135_to_check_34;

// 拆分后校验节点34传递给变量节点181的值以及对变量节点181传递过来的值
wire [5:0] value_check_34_to_variable_181;
wire enable_check_34_to_variable_181;
wire [5:0] value_variable_181_to_check_34;
wire enable_variable_181_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_181 = value_check_34_to_variable[29:24];
assign enable_check_34_to_variable_181 = enable_check_34_to_variable[4];
// 对变量节点181传递过来的值进行组合
assign value_variable_to_check_34[29:24] = value_variable_181_to_check_34;
assign enable_variable_to_check_34[4] = enable_variable_181_to_check_34;

// 拆分后校验节点34传递给变量节点229的值以及对变量节点229传递过来的值
wire [5:0] value_check_34_to_variable_229;
wire enable_check_34_to_variable_229;
wire [5:0] value_variable_229_to_check_34;
wire enable_variable_229_to_check_34;
// 对校验节点34的输出值进行拆分
assign value_check_34_to_variable_229 = value_check_34_to_variable[35:30];
assign enable_check_34_to_variable_229 = enable_check_34_to_variable[5];
// 对变量节点229传递过来的值进行组合
assign value_variable_to_check_34[35:30] = value_variable_229_to_check_34;
assign enable_variable_to_check_34[5] = enable_variable_229_to_check_34;


// 校验节点35的接口
wire [35:0] value_variable_to_check_35;
wire [35:0] value_check_35_to_variable;
wire [5:0] enable_variable_to_check_35;
wire [5:0] enable_check_35_to_variable;

// 拆分后校验节点35传递给变量节点0的值以及对变量节点0传递过来的值
wire [5:0] value_check_35_to_variable_0;
wire enable_check_35_to_variable_0;
wire [5:0] value_variable_0_to_check_35;
wire enable_variable_0_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_0 = value_check_35_to_variable[5:0];
assign enable_check_35_to_variable_0 = enable_check_35_to_variable[0];
// 对变量节点0传递过来的值进行组合
assign value_variable_to_check_35[5:0] = value_variable_0_to_check_35;
assign enable_variable_to_check_35[0] = enable_variable_0_to_check_35;

// 拆分后校验节点35传递给变量节点64的值以及对变量节点64传递过来的值
wire [5:0] value_check_35_to_variable_64;
wire enable_check_35_to_variable_64;
wire [5:0] value_variable_64_to_check_35;
wire enable_variable_64_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_64 = value_check_35_to_variable[11:6];
assign enable_check_35_to_variable_64 = enable_check_35_to_variable[1];
// 对变量节点64传递过来的值进行组合
assign value_variable_to_check_35[11:6] = value_variable_64_to_check_35;
assign enable_variable_to_check_35[1] = enable_variable_64_to_check_35;

// 拆分后校验节点35传递给变量节点113的值以及对变量节点113传递过来的值
wire [5:0] value_check_35_to_variable_113;
wire enable_check_35_to_variable_113;
wire [5:0] value_variable_113_to_check_35;
wire enable_variable_113_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_113 = value_check_35_to_variable[17:12];
assign enable_check_35_to_variable_113 = enable_check_35_to_variable[2];
// 对变量节点113传递过来的值进行组合
assign value_variable_to_check_35[17:12] = value_variable_113_to_check_35;
assign enable_variable_to_check_35[2] = enable_variable_113_to_check_35;

// 拆分后校验节点35传递给变量节点135的值以及对变量节点135传递过来的值
wire [5:0] value_check_35_to_variable_135;
wire enable_check_35_to_variable_135;
wire [5:0] value_variable_135_to_check_35;
wire enable_variable_135_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_135 = value_check_35_to_variable[23:18];
assign enable_check_35_to_variable_135 = enable_check_35_to_variable[3];
// 对变量节点135传递过来的值进行组合
assign value_variable_to_check_35[23:18] = value_variable_135_to_check_35;
assign enable_variable_to_check_35[3] = enable_variable_135_to_check_35;

// 拆分后校验节点35传递给变量节点197的值以及对变量节点197传递过来的值
wire [5:0] value_check_35_to_variable_197;
wire enable_check_35_to_variable_197;
wire [5:0] value_variable_197_to_check_35;
wire enable_variable_197_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_197 = value_check_35_to_variable[29:24];
assign enable_check_35_to_variable_197 = enable_check_35_to_variable[4];
// 对变量节点197传递过来的值进行组合
assign value_variable_to_check_35[29:24] = value_variable_197_to_check_35;
assign enable_variable_to_check_35[4] = enable_variable_197_to_check_35;

// 拆分后校验节点35传递给变量节点230的值以及对变量节点230传递过来的值
wire [5:0] value_check_35_to_variable_230;
wire enable_check_35_to_variable_230;
wire [5:0] value_variable_230_to_check_35;
wire enable_variable_230_to_check_35;
// 对校验节点35的输出值进行拆分
assign value_check_35_to_variable_230 = value_check_35_to_variable[35:30];
assign enable_check_35_to_variable_230 = enable_check_35_to_variable[5];
// 对变量节点230传递过来的值进行组合
assign value_variable_to_check_35[35:30] = value_variable_230_to_check_35;
assign enable_variable_to_check_35[5] = enable_variable_230_to_check_35;


// 校验节点36的接口
wire [35:0] value_variable_to_check_36;
wire [35:0] value_check_36_to_variable;
wire [5:0] enable_variable_to_check_36;
wire [5:0] enable_check_36_to_variable;

// 拆分后校验节点36传递给变量节点20的值以及对变量节点20传递过来的值
wire [5:0] value_check_36_to_variable_20;
wire enable_check_36_to_variable_20;
wire [5:0] value_variable_20_to_check_36;
wire enable_variable_20_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_20 = value_check_36_to_variable[5:0];
assign enable_check_36_to_variable_20 = enable_check_36_to_variable[0];
// 对变量节点20传递过来的值进行组合
assign value_variable_to_check_36[5:0] = value_variable_20_to_check_36;
assign enable_variable_to_check_36[0] = enable_variable_20_to_check_36;

// 拆分后校验节点36传递给变量节点68的值以及对变量节点68传递过来的值
wire [5:0] value_check_36_to_variable_68;
wire enable_check_36_to_variable_68;
wire [5:0] value_variable_68_to_check_36;
wire enable_variable_68_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_68 = value_check_36_to_variable[11:6];
assign enable_check_36_to_variable_68 = enable_check_36_to_variable[1];
// 对变量节点68传递过来的值进行组合
assign value_variable_to_check_36[11:6] = value_variable_68_to_check_36;
assign enable_variable_to_check_36[1] = enable_variable_68_to_check_36;

// 拆分后校验节点36传递给变量节点89的值以及对变量节点89传递过来的值
wire [5:0] value_check_36_to_variable_89;
wire enable_check_36_to_variable_89;
wire [5:0] value_variable_89_to_check_36;
wire enable_variable_89_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_89 = value_check_36_to_variable[17:12];
assign enable_check_36_to_variable_89 = enable_check_36_to_variable[2];
// 对变量节点89传递过来的值进行组合
assign value_variable_to_check_36[17:12] = value_variable_89_to_check_36;
assign enable_variable_to_check_36[2] = enable_variable_89_to_check_36;

// 拆分后校验节点36传递给变量节点138的值以及对变量节点138传递过来的值
wire [5:0] value_check_36_to_variable_138;
wire enable_check_36_to_variable_138;
wire [5:0] value_variable_138_to_check_36;
wire enable_variable_138_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_138 = value_check_36_to_variable[23:18];
assign enable_check_36_to_variable_138 = enable_check_36_to_variable[3];
// 对变量节点138传递过来的值进行组合
assign value_variable_to_check_36[23:18] = value_variable_138_to_check_36;
assign enable_variable_to_check_36[3] = enable_variable_138_to_check_36;

// 拆分后校验节点36传递给变量节点198的值以及对变量节点198传递过来的值
wire [5:0] value_check_36_to_variable_198;
wire enable_check_36_to_variable_198;
wire [5:0] value_variable_198_to_check_36;
wire enable_variable_198_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_198 = value_check_36_to_variable[29:24];
assign enable_check_36_to_variable_198 = enable_check_36_to_variable[4];
// 对变量节点198传递过来的值进行组合
assign value_variable_to_check_36[29:24] = value_variable_198_to_check_36;
assign enable_variable_to_check_36[4] = enable_variable_198_to_check_36;

// 拆分后校验节点36传递给变量节点238的值以及对变量节点238传递过来的值
wire [5:0] value_check_36_to_variable_238;
wire enable_check_36_to_variable_238;
wire [5:0] value_variable_238_to_check_36;
wire enable_variable_238_to_check_36;
// 对校验节点36的输出值进行拆分
assign value_check_36_to_variable_238 = value_check_36_to_variable[35:30];
assign enable_check_36_to_variable_238 = enable_check_36_to_variable[5];
// 对变量节点238传递过来的值进行组合
assign value_variable_to_check_36[35:30] = value_variable_238_to_check_36;
assign enable_variable_to_check_36[5] = enable_variable_238_to_check_36;


// 校验节点37的接口
wire [35:0] value_variable_to_check_37;
wire [35:0] value_check_37_to_variable;
wire [5:0] enable_variable_to_check_37;
wire [5:0] enable_check_37_to_variable;

// 拆分后校验节点37传递给变量节点19的值以及对变量节点19传递过来的值
wire [5:0] value_check_37_to_variable_19;
wire enable_check_37_to_variable_19;
wire [5:0] value_variable_19_to_check_37;
wire enable_variable_19_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_19 = value_check_37_to_variable[5:0];
assign enable_check_37_to_variable_19 = enable_check_37_to_variable[0];
// 对变量节点19传递过来的值进行组合
assign value_variable_to_check_37[5:0] = value_variable_19_to_check_37;
assign enable_variable_to_check_37[0] = enable_variable_19_to_check_37;

// 拆分后校验节点37传递给变量节点67的值以及对变量节点67传递过来的值
wire [5:0] value_check_37_to_variable_67;
wire enable_check_37_to_variable_67;
wire [5:0] value_variable_67_to_check_37;
wire enable_variable_67_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_67 = value_check_37_to_variable[11:6];
assign enable_check_37_to_variable_67 = enable_check_37_to_variable[1];
// 对变量节点67传递过来的值进行组合
assign value_variable_to_check_37[11:6] = value_variable_67_to_check_37;
assign enable_variable_to_check_37[1] = enable_variable_67_to_check_37;

// 拆分后校验节点37传递给变量节点101的值以及对变量节点101传递过来的值
wire [5:0] value_check_37_to_variable_101;
wire enable_check_37_to_variable_101;
wire [5:0] value_variable_101_to_check_37;
wire enable_variable_101_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_101 = value_check_37_to_variable[17:12];
assign enable_check_37_to_variable_101 = enable_check_37_to_variable[2];
// 对变量节点101传递过来的值进行组合
assign value_variable_to_check_37[17:12] = value_variable_101_to_check_37;
assign enable_variable_to_check_37[2] = enable_variable_101_to_check_37;

// 拆分后校验节点37传递给变量节点129的值以及对变量节点129传递过来的值
wire [5:0] value_check_37_to_variable_129;
wire enable_check_37_to_variable_129;
wire [5:0] value_variable_129_to_check_37;
wire enable_variable_129_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_129 = value_check_37_to_variable[23:18];
assign enable_check_37_to_variable_129 = enable_check_37_to_variable[3];
// 对变量节点129传递过来的值进行组合
assign value_variable_to_check_37[23:18] = value_variable_129_to_check_37;
assign enable_variable_to_check_37[3] = enable_variable_129_to_check_37;

// 拆分后校验节点37传递给变量节点189的值以及对变量节点189传递过来的值
wire [5:0] value_check_37_to_variable_189;
wire enable_check_37_to_variable_189;
wire [5:0] value_variable_189_to_check_37;
wire enable_variable_189_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_189 = value_check_37_to_variable[29:24];
assign enable_check_37_to_variable_189 = enable_check_37_to_variable[4];
// 对变量节点189传递过来的值进行组合
assign value_variable_to_check_37[29:24] = value_variable_189_to_check_37;
assign enable_variable_to_check_37[4] = enable_variable_189_to_check_37;

// 拆分后校验节点37传递给变量节点213的值以及对变量节点213传递过来的值
wire [5:0] value_check_37_to_variable_213;
wire enable_check_37_to_variable_213;
wire [5:0] value_variable_213_to_check_37;
wire enable_variable_213_to_check_37;
// 对校验节点37的输出值进行拆分
assign value_check_37_to_variable_213 = value_check_37_to_variable[35:30];
assign enable_check_37_to_variable_213 = enable_check_37_to_variable[5];
// 对变量节点213传递过来的值进行组合
assign value_variable_to_check_37[35:30] = value_variable_213_to_check_37;
assign enable_variable_to_check_37[5] = enable_variable_213_to_check_37;


// 校验节点38的接口
wire [35:0] value_variable_to_check_38;
wire [35:0] value_check_38_to_variable;
wire [5:0] enable_variable_to_check_38;
wire [5:0] enable_check_38_to_variable;

// 拆分后校验节点38传递给变量节点27的值以及对变量节点27传递过来的值
wire [5:0] value_check_38_to_variable_27;
wire enable_check_38_to_variable_27;
wire [5:0] value_variable_27_to_check_38;
wire enable_variable_27_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_27 = value_check_38_to_variable[5:0];
assign enable_check_38_to_variable_27 = enable_check_38_to_variable[0];
// 对变量节点27传递过来的值进行组合
assign value_variable_to_check_38[5:0] = value_variable_27_to_check_38;
assign enable_variable_to_check_38[0] = enable_variable_27_to_check_38;

// 拆分后校验节点38传递给变量节点69的值以及对变量节点69传递过来的值
wire [5:0] value_check_38_to_variable_69;
wire enable_check_38_to_variable_69;
wire [5:0] value_variable_69_to_check_38;
wire enable_variable_69_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_69 = value_check_38_to_variable[11:6];
assign enable_check_38_to_variable_69 = enable_check_38_to_variable[1];
// 对变量节点69传递过来的值进行组合
assign value_variable_to_check_38[11:6] = value_variable_69_to_check_38;
assign enable_variable_to_check_38[1] = enable_variable_69_to_check_38;

// 拆分后校验节点38传递给变量节点114的值以及对变量节点114传递过来的值
wire [5:0] value_check_38_to_variable_114;
wire enable_check_38_to_variable_114;
wire [5:0] value_variable_114_to_check_38;
wire enable_variable_114_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_114 = value_check_38_to_variable[17:12];
assign enable_check_38_to_variable_114 = enable_check_38_to_variable[2];
// 对变量节点114传递过来的值进行组合
assign value_variable_to_check_38[17:12] = value_variable_114_to_check_38;
assign enable_variable_to_check_38[2] = enable_variable_114_to_check_38;

// 拆分后校验节点38传递给变量节点155的值以及对变量节点155传递过来的值
wire [5:0] value_check_38_to_variable_155;
wire enable_check_38_to_variable_155;
wire [5:0] value_variable_155_to_check_38;
wire enable_variable_155_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_155 = value_check_38_to_variable[23:18];
assign enable_check_38_to_variable_155 = enable_check_38_to_variable[3];
// 对变量节点155传递过来的值进行组合
assign value_variable_to_check_38[23:18] = value_variable_155_to_check_38;
assign enable_variable_to_check_38[3] = enable_variable_155_to_check_38;

// 拆分后校验节点38传递给变量节点172的值以及对变量节点172传递过来的值
wire [5:0] value_check_38_to_variable_172;
wire enable_check_38_to_variable_172;
wire [5:0] value_variable_172_to_check_38;
wire enable_variable_172_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_172 = value_check_38_to_variable[29:24];
assign enable_check_38_to_variable_172 = enable_check_38_to_variable[4];
// 对变量节点172传递过来的值进行组合
assign value_variable_to_check_38[29:24] = value_variable_172_to_check_38;
assign enable_variable_to_check_38[4] = enable_variable_172_to_check_38;

// 拆分后校验节点38传递给变量节点221的值以及对变量节点221传递过来的值
wire [5:0] value_check_38_to_variable_221;
wire enable_check_38_to_variable_221;
wire [5:0] value_variable_221_to_check_38;
wire enable_variable_221_to_check_38;
// 对校验节点38的输出值进行拆分
assign value_check_38_to_variable_221 = value_check_38_to_variable[35:30];
assign enable_check_38_to_variable_221 = enable_check_38_to_variable[5];
// 对变量节点221传递过来的值进行组合
assign value_variable_to_check_38[35:30] = value_variable_221_to_check_38;
assign enable_variable_to_check_38[5] = enable_variable_221_to_check_38;


// 校验节点39的接口
wire [35:0] value_variable_to_check_39;
wire [35:0] value_check_39_to_variable;
wire [5:0] enable_variable_to_check_39;
wire [5:0] enable_check_39_to_variable;

// 拆分后校验节点39传递给变量节点21的值以及对变量节点21传递过来的值
wire [5:0] value_check_39_to_variable_21;
wire enable_check_39_to_variable_21;
wire [5:0] value_variable_21_to_check_39;
wire enable_variable_21_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_21 = value_check_39_to_variable[5:0];
assign enable_check_39_to_variable_21 = enable_check_39_to_variable[0];
// 对变量节点21传递过来的值进行组合
assign value_variable_to_check_39[5:0] = value_variable_21_to_check_39;
assign enable_variable_to_check_39[0] = enable_variable_21_to_check_39;

// 拆分后校验节点39传递给变量节点70的值以及对变量节点70传递过来的值
wire [5:0] value_check_39_to_variable_70;
wire enable_check_39_to_variable_70;
wire [5:0] value_variable_70_to_check_39;
wire enable_variable_70_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_70 = value_check_39_to_variable[11:6];
assign enable_check_39_to_variable_70 = enable_check_39_to_variable[1];
// 对变量节点70传递过来的值进行组合
assign value_variable_to_check_39[11:6] = value_variable_70_to_check_39;
assign enable_variable_to_check_39[1] = enable_variable_70_to_check_39;

// 拆分后校验节点39传递给变量节点115的值以及对变量节点115传递过来的值
wire [5:0] value_check_39_to_variable_115;
wire enable_check_39_to_variable_115;
wire [5:0] value_variable_115_to_check_39;
wire enable_variable_115_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_115 = value_check_39_to_variable[17:12];
assign enable_check_39_to_variable_115 = enable_check_39_to_variable[2];
// 对变量节点115传递过来的值进行组合
assign value_variable_to_check_39[17:12] = value_variable_115_to_check_39;
assign enable_variable_to_check_39[2] = enable_variable_115_to_check_39;

// 拆分后校验节点39传递给变量节点146的值以及对变量节点146传递过来的值
wire [5:0] value_check_39_to_variable_146;
wire enable_check_39_to_variable_146;
wire [5:0] value_variable_146_to_check_39;
wire enable_variable_146_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_146 = value_check_39_to_variable[23:18];
assign enable_check_39_to_variable_146 = enable_check_39_to_variable[3];
// 对变量节点146传递过来的值进行组合
assign value_variable_to_check_39[23:18] = value_variable_146_to_check_39;
assign enable_variable_to_check_39[3] = enable_variable_146_to_check_39;

// 拆分后校验节点39传递给变量节点199的值以及对变量节点199传递过来的值
wire [5:0] value_check_39_to_variable_199;
wire enable_check_39_to_variable_199;
wire [5:0] value_variable_199_to_check_39;
wire enable_variable_199_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_199 = value_check_39_to_variable[29:24];
assign enable_check_39_to_variable_199 = enable_check_39_to_variable[4];
// 对变量节点199传递过来的值进行组合
assign value_variable_to_check_39[29:24] = value_variable_199_to_check_39;
assign enable_variable_to_check_39[4] = enable_variable_199_to_check_39;

// 拆分后校验节点39传递给变量节点239的值以及对变量节点239传递过来的值
wire [5:0] value_check_39_to_variable_239;
wire enable_check_39_to_variable_239;
wire [5:0] value_variable_239_to_check_39;
wire enable_variable_239_to_check_39;
// 对校验节点39的输出值进行拆分
assign value_check_39_to_variable_239 = value_check_39_to_variable[35:30];
assign enable_check_39_to_variable_239 = enable_check_39_to_variable[5];
// 对变量节点239传递过来的值进行组合
assign value_variable_to_check_39[35:30] = value_variable_239_to_check_39;
assign enable_variable_to_check_39[5] = enable_variable_239_to_check_39;


// 校验节点40的接口
wire [35:0] value_variable_to_check_40;
wire [35:0] value_check_40_to_variable;
wire [5:0] enable_variable_to_check_40;
wire [5:0] enable_check_40_to_variable;

// 拆分后校验节点40传递给变量节点15的值以及对变量节点15传递过来的值
wire [5:0] value_check_40_to_variable_15;
wire enable_check_40_to_variable_15;
wire [5:0] value_variable_15_to_check_40;
wire enable_variable_15_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_15 = value_check_40_to_variable[5:0];
assign enable_check_40_to_variable_15 = enable_check_40_to_variable[0];
// 对变量节点15传递过来的值进行组合
assign value_variable_to_check_40[5:0] = value_variable_15_to_check_40;
assign enable_variable_to_check_40[0] = enable_variable_15_to_check_40;

// 拆分后校验节点40传递给变量节点71的值以及对变量节点71传递过来的值
wire [5:0] value_check_40_to_variable_71;
wire enable_check_40_to_variable_71;
wire [5:0] value_variable_71_to_check_40;
wire enable_variable_71_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_71 = value_check_40_to_variable[11:6];
assign enable_check_40_to_variable_71 = enable_check_40_to_variable[1];
// 对变量节点71传递过来的值进行组合
assign value_variable_to_check_40[11:6] = value_variable_71_to_check_40;
assign enable_variable_to_check_40[1] = enable_variable_71_to_check_40;

// 拆分后校验节点40传递给变量节点116的值以及对变量节点116传递过来的值
wire [5:0] value_check_40_to_variable_116;
wire enable_check_40_to_variable_116;
wire [5:0] value_variable_116_to_check_40;
wire enable_variable_116_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_116 = value_check_40_to_variable[17:12];
assign enable_check_40_to_variable_116 = enable_check_40_to_variable[2];
// 对变量节点116传递过来的值进行组合
assign value_variable_to_check_40[17:12] = value_variable_116_to_check_40;
assign enable_variable_to_check_40[2] = enable_variable_116_to_check_40;

// 拆分后校验节点40传递给变量节点139的值以及对变量节点139传递过来的值
wire [5:0] value_check_40_to_variable_139;
wire enable_check_40_to_variable_139;
wire [5:0] value_variable_139_to_check_40;
wire enable_variable_139_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_139 = value_check_40_to_variable[23:18];
assign enable_check_40_to_variable_139 = enable_check_40_to_variable[3];
// 对变量节点139传递过来的值进行组合
assign value_variable_to_check_40[23:18] = value_variable_139_to_check_40;
assign enable_variable_to_check_40[3] = enable_variable_139_to_check_40;

// 拆分后校验节点40传递给变量节点200的值以及对变量节点200传递过来的值
wire [5:0] value_check_40_to_variable_200;
wire enable_check_40_to_variable_200;
wire [5:0] value_variable_200_to_check_40;
wire enable_variable_200_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_200 = value_check_40_to_variable[29:24];
assign enable_check_40_to_variable_200 = enable_check_40_to_variable[4];
// 对变量节点200传递过来的值进行组合
assign value_variable_to_check_40[29:24] = value_variable_200_to_check_40;
assign enable_variable_to_check_40[4] = enable_variable_200_to_check_40;

// 拆分后校验节点40传递给变量节点240的值以及对变量节点240传递过来的值
wire [5:0] value_check_40_to_variable_240;
wire enable_check_40_to_variable_240;
wire [5:0] value_variable_240_to_check_40;
wire enable_variable_240_to_check_40;
// 对校验节点40的输出值进行拆分
assign value_check_40_to_variable_240 = value_check_40_to_variable[35:30];
assign enable_check_40_to_variable_240 = enable_check_40_to_variable[5];
// 对变量节点240传递过来的值进行组合
assign value_variable_to_check_40[35:30] = value_variable_240_to_check_40;
assign enable_variable_to_check_40[5] = enable_variable_240_to_check_40;


// 校验节点41的接口
wire [35:0] value_variable_to_check_41;
wire [35:0] value_check_41_to_variable;
wire [5:0] enable_variable_to_check_41;
wire [5:0] enable_check_41_to_variable;

// 拆分后校验节点41传递给变量节点20的值以及对变量节点20传递过来的值
wire [5:0] value_check_41_to_variable_20;
wire enable_check_41_to_variable_20;
wire [5:0] value_variable_20_to_check_41;
wire enable_variable_20_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_20 = value_check_41_to_variable[5:0];
assign enable_check_41_to_variable_20 = enable_check_41_to_variable[0];
// 对变量节点20传递过来的值进行组合
assign value_variable_to_check_41[5:0] = value_variable_20_to_check_41;
assign enable_variable_to_check_41[0] = enable_variable_20_to_check_41;

// 拆分后校验节点41传递给变量节点64的值以及对变量节点64传递过来的值
wire [5:0] value_check_41_to_variable_64;
wire enable_check_41_to_variable_64;
wire [5:0] value_variable_64_to_check_41;
wire enable_variable_64_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_64 = value_check_41_to_variable[11:6];
assign enable_check_41_to_variable_64 = enable_check_41_to_variable[1];
// 对变量节点64传递过来的值进行组合
assign value_variable_to_check_41[11:6] = value_variable_64_to_check_41;
assign enable_variable_to_check_41[1] = enable_variable_64_to_check_41;

// 拆分后校验节点41传递给变量节点90的值以及对变量节点90传递过来的值
wire [5:0] value_check_41_to_variable_90;
wire enable_check_41_to_variable_90;
wire [5:0] value_variable_90_to_check_41;
wire enable_variable_90_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_90 = value_check_41_to_variable[17:12];
assign enable_check_41_to_variable_90 = enable_check_41_to_variable[2];
// 对变量节点90传递过来的值进行组合
assign value_variable_to_check_41[17:12] = value_variable_90_to_check_41;
assign enable_variable_to_check_41[2] = enable_variable_90_to_check_41;

// 拆分后校验节点41传递给变量节点142的值以及对变量节点142传递过来的值
wire [5:0] value_check_41_to_variable_142;
wire enable_check_41_to_variable_142;
wire [5:0] value_variable_142_to_check_41;
wire enable_variable_142_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_142 = value_check_41_to_variable[23:18];
assign enable_check_41_to_variable_142 = enable_check_41_to_variable[3];
// 对变量节点142传递过来的值进行组合
assign value_variable_to_check_41[23:18] = value_variable_142_to_check_41;
assign enable_variable_to_check_41[3] = enable_variable_142_to_check_41;

// 拆分后校验节点41传递给变量节点201的值以及对变量节点201传递过来的值
wire [5:0] value_check_41_to_variable_201;
wire enable_check_41_to_variable_201;
wire [5:0] value_variable_201_to_check_41;
wire enable_variable_201_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_201 = value_check_41_to_variable[29:24];
assign enable_check_41_to_variable_201 = enable_check_41_to_variable[4];
// 对变量节点201传递过来的值进行组合
assign value_variable_to_check_41[29:24] = value_variable_201_to_check_41;
assign enable_variable_to_check_41[4] = enable_variable_201_to_check_41;

// 拆分后校验节点41传递给变量节点241的值以及对变量节点241传递过来的值
wire [5:0] value_check_41_to_variable_241;
wire enable_check_41_to_variable_241;
wire [5:0] value_variable_241_to_check_41;
wire enable_variable_241_to_check_41;
// 对校验节点41的输出值进行拆分
assign value_check_41_to_variable_241 = value_check_41_to_variable[35:30];
assign enable_check_41_to_variable_241 = enable_check_41_to_variable[5];
// 对变量节点241传递过来的值进行组合
assign value_variable_to_check_41[35:30] = value_variable_241_to_check_41;
assign enable_variable_to_check_41[5] = enable_variable_241_to_check_41;


// 校验节点42的接口
wire [35:0] value_variable_to_check_42;
wire [35:0] value_check_42_to_variable;
wire [5:0] enable_variable_to_check_42;
wire [5:0] enable_check_42_to_variable;

// 拆分后校验节点42传递给变量节点28的值以及对变量节点28传递过来的值
wire [5:0] value_check_42_to_variable_28;
wire enable_check_42_to_variable_28;
wire [5:0] value_variable_28_to_check_42;
wire enable_variable_28_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_28 = value_check_42_to_variable[5:0];
assign enable_check_42_to_variable_28 = enable_check_42_to_variable[0];
// 对变量节点28传递过来的值进行组合
assign value_variable_to_check_42[5:0] = value_variable_28_to_check_42;
assign enable_variable_to_check_42[0] = enable_variable_28_to_check_42;

// 拆分后校验节点42传递给变量节点72的值以及对变量节点72传递过来的值
wire [5:0] value_check_42_to_variable_72;
wire enable_check_42_to_variable_72;
wire [5:0] value_variable_72_to_check_42;
wire enable_variable_72_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_72 = value_check_42_to_variable[11:6];
assign enable_check_42_to_variable_72 = enable_check_42_to_variable[1];
// 对变量节点72传递过来的值进行组合
assign value_variable_to_check_42[11:6] = value_variable_72_to_check_42;
assign enable_variable_to_check_42[1] = enable_variable_72_to_check_42;

// 拆分后校验节点42传递给变量节点92的值以及对变量节点92传递过来的值
wire [5:0] value_check_42_to_variable_92;
wire enable_check_42_to_variable_92;
wire [5:0] value_variable_92_to_check_42;
wire enable_variable_92_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_92 = value_check_42_to_variable[17:12];
assign enable_check_42_to_variable_92 = enable_check_42_to_variable[2];
// 对变量节点92传递过来的值进行组合
assign value_variable_to_check_42[17:12] = value_variable_92_to_check_42;
assign enable_variable_to_check_42[2] = enable_variable_92_to_check_42;

// 拆分后校验节点42传递给变量节点144的值以及对变量节点144传递过来的值
wire [5:0] value_check_42_to_variable_144;
wire enable_check_42_to_variable_144;
wire [5:0] value_variable_144_to_check_42;
wire enable_variable_144_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_144 = value_check_42_to_variable[23:18];
assign enable_check_42_to_variable_144 = enable_check_42_to_variable[3];
// 对变量节点144传递过来的值进行组合
assign value_variable_to_check_42[23:18] = value_variable_144_to_check_42;
assign enable_variable_to_check_42[3] = enable_variable_144_to_check_42;

// 拆分后校验节点42传递给变量节点202的值以及对变量节点202传递过来的值
wire [5:0] value_check_42_to_variable_202;
wire enable_check_42_to_variable_202;
wire [5:0] value_variable_202_to_check_42;
wire enable_variable_202_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_202 = value_check_42_to_variable[29:24];
assign enable_check_42_to_variable_202 = enable_check_42_to_variable[4];
// 对变量节点202传递过来的值进行组合
assign value_variable_to_check_42[29:24] = value_variable_202_to_check_42;
assign enable_variable_to_check_42[4] = enable_variable_202_to_check_42;

// 拆分后校验节点42传递给变量节点232的值以及对变量节点232传递过来的值
wire [5:0] value_check_42_to_variable_232;
wire enable_check_42_to_variable_232;
wire [5:0] value_variable_232_to_check_42;
wire enable_variable_232_to_check_42;
// 对校验节点42的输出值进行拆分
assign value_check_42_to_variable_232 = value_check_42_to_variable[35:30];
assign enable_check_42_to_variable_232 = enable_check_42_to_variable[5];
// 对变量节点232传递过来的值进行组合
assign value_variable_to_check_42[35:30] = value_variable_232_to_check_42;
assign enable_variable_to_check_42[5] = enable_variable_232_to_check_42;


// 校验节点43的接口
wire [35:0] value_variable_to_check_43;
wire [35:0] value_check_43_to_variable;
wire [5:0] enable_variable_to_check_43;
wire [5:0] enable_check_43_to_variable;

// 拆分后校验节点43传递给变量节点29的值以及对变量节点29传递过来的值
wire [5:0] value_check_43_to_variable_29;
wire enable_check_43_to_variable_29;
wire [5:0] value_variable_29_to_check_43;
wire enable_variable_29_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_29 = value_check_43_to_variable[5:0];
assign enable_check_43_to_variable_29 = enable_check_43_to_variable[0];
// 对变量节点29传递过来的值进行组合
assign value_variable_to_check_43[5:0] = value_variable_29_to_check_43;
assign enable_variable_to_check_43[0] = enable_variable_29_to_check_43;

// 拆分后校验节点43传递给变量节点73的值以及对变量节点73传递过来的值
wire [5:0] value_check_43_to_variable_73;
wire enable_check_43_to_variable_73;
wire [5:0] value_variable_73_to_check_43;
wire enable_variable_73_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_73 = value_check_43_to_variable[11:6];
assign enable_check_43_to_variable_73 = enable_check_43_to_variable[1];
// 对变量节点73传递过来的值进行组合
assign value_variable_to_check_43[11:6] = value_variable_73_to_check_43;
assign enable_variable_to_check_43[1] = enable_variable_73_to_check_43;

// 拆分后校验节点43传递给变量节点117的值以及对变量节点117传递过来的值
wire [5:0] value_check_43_to_variable_117;
wire enable_check_43_to_variable_117;
wire [5:0] value_variable_117_to_check_43;
wire enable_variable_117_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_117 = value_check_43_to_variable[17:12];
assign enable_check_43_to_variable_117 = enable_check_43_to_variable[2];
// 对变量节点117传递过来的值进行组合
assign value_variable_to_check_43[17:12] = value_variable_117_to_check_43;
assign enable_variable_to_check_43[2] = enable_variable_117_to_check_43;

// 拆分后校验节点43传递给变量节点143的值以及对变量节点143传递过来的值
wire [5:0] value_check_43_to_variable_143;
wire enable_check_43_to_variable_143;
wire [5:0] value_variable_143_to_check_43;
wire enable_variable_143_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_143 = value_check_43_to_variable[23:18];
assign enable_check_43_to_variable_143 = enable_check_43_to_variable[3];
// 对变量节点143传递过来的值进行组合
assign value_variable_to_check_43[23:18] = value_variable_143_to_check_43;
assign enable_variable_to_check_43[3] = enable_variable_143_to_check_43;

// 拆分后校验节点43传递给变量节点176的值以及对变量节点176传递过来的值
wire [5:0] value_check_43_to_variable_176;
wire enable_check_43_to_variable_176;
wire [5:0] value_variable_176_to_check_43;
wire enable_variable_176_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_176 = value_check_43_to_variable[29:24];
assign enable_check_43_to_variable_176 = enable_check_43_to_variable[4];
// 对变量节点176传递过来的值进行组合
assign value_variable_to_check_43[29:24] = value_variable_176_to_check_43;
assign enable_variable_to_check_43[4] = enable_variable_176_to_check_43;

// 拆分后校验节点43传递给变量节点219的值以及对变量节点219传递过来的值
wire [5:0] value_check_43_to_variable_219;
wire enable_check_43_to_variable_219;
wire [5:0] value_variable_219_to_check_43;
wire enable_variable_219_to_check_43;
// 对校验节点43的输出值进行拆分
assign value_check_43_to_variable_219 = value_check_43_to_variable[35:30];
assign enable_check_43_to_variable_219 = enable_check_43_to_variable[5];
// 对变量节点219传递过来的值进行组合
assign value_variable_to_check_43[35:30] = value_variable_219_to_check_43;
assign enable_variable_to_check_43[5] = enable_variable_219_to_check_43;


// 校验节点44的接口
wire [35:0] value_variable_to_check_44;
wire [35:0] value_check_44_to_variable;
wire [5:0] enable_variable_to_check_44;
wire [5:0] enable_check_44_to_variable;

// 拆分后校验节点44传递给变量节点2的值以及对变量节点2传递过来的值
wire [5:0] value_check_44_to_variable_2;
wire enable_check_44_to_variable_2;
wire [5:0] value_variable_2_to_check_44;
wire enable_variable_2_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_2 = value_check_44_to_variable[5:0];
assign enable_check_44_to_variable_2 = enable_check_44_to_variable[0];
// 对变量节点2传递过来的值进行组合
assign value_variable_to_check_44[5:0] = value_variable_2_to_check_44;
assign enable_variable_to_check_44[0] = enable_variable_2_to_check_44;

// 拆分后校验节点44传递给变量节点66的值以及对变量节点66传递过来的值
wire [5:0] value_check_44_to_variable_66;
wire enable_check_44_to_variable_66;
wire [5:0] value_variable_66_to_check_44;
wire enable_variable_66_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_66 = value_check_44_to_variable[11:6];
assign enable_check_44_to_variable_66 = enable_check_44_to_variable[1];
// 对变量节点66传递过来的值进行组合
assign value_variable_to_check_44[11:6] = value_variable_66_to_check_44;
assign enable_variable_to_check_44[1] = enable_variable_66_to_check_44;

// 拆分后校验节点44传递给变量节点106的值以及对变量节点106传递过来的值
wire [5:0] value_check_44_to_variable_106;
wire enable_check_44_to_variable_106;
wire [5:0] value_variable_106_to_check_44;
wire enable_variable_106_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_106 = value_check_44_to_variable[17:12];
assign enable_check_44_to_variable_106 = enable_check_44_to_variable[2];
// 对变量节点106传递过来的值进行组合
assign value_variable_to_check_44[17:12] = value_variable_106_to_check_44;
assign enable_variable_to_check_44[2] = enable_variable_106_to_check_44;

// 拆分后校验节点44传递给变量节点157的值以及对变量节点157传递过来的值
wire [5:0] value_check_44_to_variable_157;
wire enable_check_44_to_variable_157;
wire [5:0] value_variable_157_to_check_44;
wire enable_variable_157_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_157 = value_check_44_to_variable[23:18];
assign enable_check_44_to_variable_157 = enable_check_44_to_variable[3];
// 对变量节点157传递过来的值进行组合
assign value_variable_to_check_44[23:18] = value_variable_157_to_check_44;
assign enable_variable_to_check_44[3] = enable_variable_157_to_check_44;

// 拆分后校验节点44传递给变量节点203的值以及对变量节点203传递过来的值
wire [5:0] value_check_44_to_variable_203;
wire enable_check_44_to_variable_203;
wire [5:0] value_variable_203_to_check_44;
wire enable_variable_203_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_203 = value_check_44_to_variable[29:24];
assign enable_check_44_to_variable_203 = enable_check_44_to_variable[4];
// 对变量节点203传递过来的值进行组合
assign value_variable_to_check_44[29:24] = value_variable_203_to_check_44;
assign enable_variable_to_check_44[4] = enable_variable_203_to_check_44;

// 拆分后校验节点44传递给变量节点231的值以及对变量节点231传递过来的值
wire [5:0] value_check_44_to_variable_231;
wire enable_check_44_to_variable_231;
wire [5:0] value_variable_231_to_check_44;
wire enable_variable_231_to_check_44;
// 对校验节点44的输出值进行拆分
assign value_check_44_to_variable_231 = value_check_44_to_variable[35:30];
assign enable_check_44_to_variable_231 = enable_check_44_to_variable[5];
// 对变量节点231传递过来的值进行组合
assign value_variable_to_check_44[35:30] = value_variable_231_to_check_44;
assign enable_variable_to_check_44[5] = enable_variable_231_to_check_44;


// 校验节点45的接口
wire [35:0] value_variable_to_check_45;
wire [35:0] value_check_45_to_variable;
wire [5:0] enable_variable_to_check_45;
wire [5:0] enable_check_45_to_variable;

// 拆分后校验节点45传递给变量节点30的值以及对变量节点30传递过来的值
wire [5:0] value_check_45_to_variable_30;
wire enable_check_45_to_variable_30;
wire [5:0] value_variable_30_to_check_45;
wire enable_variable_30_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_30 = value_check_45_to_variable[5:0];
assign enable_check_45_to_variable_30 = enable_check_45_to_variable[0];
// 对变量节点30传递过来的值进行组合
assign value_variable_to_check_45[5:0] = value_variable_30_to_check_45;
assign enable_variable_to_check_45[0] = enable_variable_30_to_check_45;

// 拆分后校验节点45传递给变量节点62的值以及对变量节点62传递过来的值
wire [5:0] value_check_45_to_variable_62;
wire enable_check_45_to_variable_62;
wire [5:0] value_variable_62_to_check_45;
wire enable_variable_62_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_62 = value_check_45_to_variable[11:6];
assign enable_check_45_to_variable_62 = enable_check_45_to_variable[1];
// 对变量节点62传递过来的值进行组合
assign value_variable_to_check_45[11:6] = value_variable_62_to_check_45;
assign enable_variable_to_check_45[1] = enable_variable_62_to_check_45;

// 拆分后校验节点45传递给变量节点118的值以及对变量节点118传递过来的值
wire [5:0] value_check_45_to_variable_118;
wire enable_check_45_to_variable_118;
wire [5:0] value_variable_118_to_check_45;
wire enable_variable_118_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_118 = value_check_45_to_variable[17:12];
assign enable_check_45_to_variable_118 = enable_check_45_to_variable[2];
// 对变量节点118传递过来的值进行组合
assign value_variable_to_check_45[17:12] = value_variable_118_to_check_45;
assign enable_variable_to_check_45[2] = enable_variable_118_to_check_45;

// 拆分后校验节点45传递给变量节点159的值以及对变量节点159传递过来的值
wire [5:0] value_check_45_to_variable_159;
wire enable_check_45_to_variable_159;
wire [5:0] value_variable_159_to_check_45;
wire enable_variable_159_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_159 = value_check_45_to_variable[23:18];
assign enable_check_45_to_variable_159 = enable_check_45_to_variable[3];
// 对变量节点159传递过来的值进行组合
assign value_variable_to_check_45[23:18] = value_variable_159_to_check_45;
assign enable_variable_to_check_45[3] = enable_variable_159_to_check_45;

// 拆分后校验节点45传递给变量节点195的值以及对变量节点195传递过来的值
wire [5:0] value_check_45_to_variable_195;
wire enable_check_45_to_variable_195;
wire [5:0] value_variable_195_to_check_45;
wire enable_variable_195_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_195 = value_check_45_to_variable[29:24];
assign enable_check_45_to_variable_195 = enable_check_45_to_variable[4];
// 对变量节点195传递过来的值进行组合
assign value_variable_to_check_45[29:24] = value_variable_195_to_check_45;
assign enable_variable_to_check_45[4] = enable_variable_195_to_check_45;

// 拆分后校验节点45传递给变量节点227的值以及对变量节点227传递过来的值
wire [5:0] value_check_45_to_variable_227;
wire enable_check_45_to_variable_227;
wire [5:0] value_variable_227_to_check_45;
wire enable_variable_227_to_check_45;
// 对校验节点45的输出值进行拆分
assign value_check_45_to_variable_227 = value_check_45_to_variable[35:30];
assign enable_check_45_to_variable_227 = enable_check_45_to_variable[5];
// 对变量节点227传递过来的值进行组合
assign value_variable_to_check_45[35:30] = value_variable_227_to_check_45;
assign enable_variable_to_check_45[5] = enable_variable_227_to_check_45;


// 校验节点46的接口
wire [35:0] value_variable_to_check_46;
wire [35:0] value_check_46_to_variable;
wire [5:0] enable_variable_to_check_46;
wire [5:0] enable_check_46_to_variable;

// 拆分后校验节点46传递给变量节点5的值以及对变量节点5传递过来的值
wire [5:0] value_check_46_to_variable_5;
wire enable_check_46_to_variable_5;
wire [5:0] value_variable_5_to_check_46;
wire enable_variable_5_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_5 = value_check_46_to_variable[5:0];
assign enable_check_46_to_variable_5 = enable_check_46_to_variable[0];
// 对变量节点5传递过来的值进行组合
assign value_variable_to_check_46[5:0] = value_variable_5_to_check_46;
assign enable_variable_to_check_46[0] = enable_variable_5_to_check_46;

// 拆分后校验节点46传递给变量节点56的值以及对变量节点56传递过来的值
wire [5:0] value_check_46_to_variable_56;
wire enable_check_46_to_variable_56;
wire [5:0] value_variable_56_to_check_46;
wire enable_variable_56_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_56 = value_check_46_to_variable[11:6];
assign enable_check_46_to_variable_56 = enable_check_46_to_variable[1];
// 对变量节点56传递过来的值进行组合
assign value_variable_to_check_46[11:6] = value_variable_56_to_check_46;
assign enable_variable_to_check_46[1] = enable_variable_56_to_check_46;

// 拆分后校验节点46传递给变量节点87的值以及对变量节点87传递过来的值
wire [5:0] value_check_46_to_variable_87;
wire enable_check_46_to_variable_87;
wire [5:0] value_variable_87_to_check_46;
wire enable_variable_87_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_87 = value_check_46_to_variable[17:12];
assign enable_check_46_to_variable_87 = enable_check_46_to_variable[2];
// 对变量节点87传递过来的值进行组合
assign value_variable_to_check_46[17:12] = value_variable_87_to_check_46;
assign enable_variable_to_check_46[2] = enable_variable_87_to_check_46;

// 拆分后校验节点46传递给变量节点153的值以及对变量节点153传递过来的值
wire [5:0] value_check_46_to_variable_153;
wire enable_check_46_to_variable_153;
wire [5:0] value_variable_153_to_check_46;
wire enable_variable_153_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_153 = value_check_46_to_variable[23:18];
assign enable_check_46_to_variable_153 = enable_check_46_to_variable[3];
// 对变量节点153传递过来的值进行组合
assign value_variable_to_check_46[23:18] = value_variable_153_to_check_46;
assign enable_variable_to_check_46[3] = enable_variable_153_to_check_46;

// 拆分后校验节点46传递给变量节点204的值以及对变量节点204传递过来的值
wire [5:0] value_check_46_to_variable_204;
wire enable_check_46_to_variable_204;
wire [5:0] value_variable_204_to_check_46;
wire enable_variable_204_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_204 = value_check_46_to_variable[29:24];
assign enable_check_46_to_variable_204 = enable_check_46_to_variable[4];
// 对变量节点204传递过来的值进行组合
assign value_variable_to_check_46[29:24] = value_variable_204_to_check_46;
assign enable_variable_to_check_46[4] = enable_variable_204_to_check_46;

// 拆分后校验节点46传递给变量节点242的值以及对变量节点242传递过来的值
wire [5:0] value_check_46_to_variable_242;
wire enable_check_46_to_variable_242;
wire [5:0] value_variable_242_to_check_46;
wire enable_variable_242_to_check_46;
// 对校验节点46的输出值进行拆分
assign value_check_46_to_variable_242 = value_check_46_to_variable[35:30];
assign enable_check_46_to_variable_242 = enable_check_46_to_variable[5];
// 对变量节点242传递过来的值进行组合
assign value_variable_to_check_46[35:30] = value_variable_242_to_check_46;
assign enable_variable_to_check_46[5] = enable_variable_242_to_check_46;


// 校验节点47的接口
wire [35:0] value_variable_to_check_47;
wire [35:0] value_check_47_to_variable;
wire [5:0] enable_variable_to_check_47;
wire [5:0] enable_check_47_to_variable;

// 拆分后校验节点47传递给变量节点31的值以及对变量节点31传递过来的值
wire [5:0] value_check_47_to_variable_31;
wire enable_check_47_to_variable_31;
wire [5:0] value_variable_31_to_check_47;
wire enable_variable_31_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_31 = value_check_47_to_variable[5:0];
assign enable_check_47_to_variable_31 = enable_check_47_to_variable[0];
// 对变量节点31传递过来的值进行组合
assign value_variable_to_check_47[5:0] = value_variable_31_to_check_47;
assign enable_variable_to_check_47[0] = enable_variable_31_to_check_47;

// 拆分后校验节点47传递给变量节点51的值以及对变量节点51传递过来的值
wire [5:0] value_check_47_to_variable_51;
wire enable_check_47_to_variable_51;
wire [5:0] value_variable_51_to_check_47;
wire enable_variable_51_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_51 = value_check_47_to_variable[11:6];
assign enable_check_47_to_variable_51 = enable_check_47_to_variable[1];
// 对变量节点51传递过来的值进行组合
assign value_variable_to_check_47[11:6] = value_variable_51_to_check_47;
assign enable_variable_to_check_47[1] = enable_variable_51_to_check_47;

// 拆分后校验节点47传递给变量节点119的值以及对变量节点119传递过来的值
wire [5:0] value_check_47_to_variable_119;
wire enable_check_47_to_variable_119;
wire [5:0] value_variable_119_to_check_47;
wire enable_variable_119_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_119 = value_check_47_to_variable[17:12];
assign enable_check_47_to_variable_119 = enable_check_47_to_variable[2];
// 对变量节点119传递过来的值进行组合
assign value_variable_to_check_47[17:12] = value_variable_119_to_check_47;
assign enable_variable_to_check_47[2] = enable_variable_119_to_check_47;

// 拆分后校验节点47传递给变量节点143的值以及对变量节点143传递过来的值
wire [5:0] value_check_47_to_variable_143;
wire enable_check_47_to_variable_143;
wire [5:0] value_variable_143_to_check_47;
wire enable_variable_143_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_143 = value_check_47_to_variable[23:18];
assign enable_check_47_to_variable_143 = enable_check_47_to_variable[3];
// 对变量节点143传递过来的值进行组合
assign value_variable_to_check_47[23:18] = value_variable_143_to_check_47;
assign enable_variable_to_check_47[3] = enable_variable_143_to_check_47;

// 拆分后校验节点47传递给变量节点198的值以及对变量节点198传递过来的值
wire [5:0] value_check_47_to_variable_198;
wire enable_check_47_to_variable_198;
wire [5:0] value_variable_198_to_check_47;
wire enable_variable_198_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_198 = value_check_47_to_variable[29:24];
assign enable_check_47_to_variable_198 = enable_check_47_to_variable[4];
// 对变量节点198传递过来的值进行组合
assign value_variable_to_check_47[29:24] = value_variable_198_to_check_47;
assign enable_variable_to_check_47[4] = enable_variable_198_to_check_47;

// 拆分后校验节点47传递给变量节点228的值以及对变量节点228传递过来的值
wire [5:0] value_check_47_to_variable_228;
wire enable_check_47_to_variable_228;
wire [5:0] value_variable_228_to_check_47;
wire enable_variable_228_to_check_47;
// 对校验节点47的输出值进行拆分
assign value_check_47_to_variable_228 = value_check_47_to_variable[35:30];
assign enable_check_47_to_variable_228 = enable_check_47_to_variable[5];
// 对变量节点228传递过来的值进行组合
assign value_variable_to_check_47[35:30] = value_variable_228_to_check_47;
assign enable_variable_to_check_47[5] = enable_variable_228_to_check_47;


// 校验节点48的接口
wire [35:0] value_variable_to_check_48;
wire [35:0] value_check_48_to_variable;
wire [5:0] enable_variable_to_check_48;
wire [5:0] enable_check_48_to_variable;

// 拆分后校验节点48传递给变量节点21的值以及对变量节点21传递过来的值
wire [5:0] value_check_48_to_variable_21;
wire enable_check_48_to_variable_21;
wire [5:0] value_variable_21_to_check_48;
wire enable_variable_21_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_21 = value_check_48_to_variable[5:0];
assign enable_check_48_to_variable_21 = enable_check_48_to_variable[0];
// 对变量节点21传递过来的值进行组合
assign value_variable_to_check_48[5:0] = value_variable_21_to_check_48;
assign enable_variable_to_check_48[0] = enable_variable_21_to_check_48;

// 拆分后校验节点48传递给变量节点46的值以及对变量节点46传递过来的值
wire [5:0] value_check_48_to_variable_46;
wire enable_check_48_to_variable_46;
wire [5:0] value_variable_46_to_check_48;
wire enable_variable_46_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_46 = value_check_48_to_variable[11:6];
assign enable_check_48_to_variable_46 = enable_check_48_to_variable[1];
// 对变量节点46传递过来的值进行组合
assign value_variable_to_check_48[11:6] = value_variable_46_to_check_48;
assign enable_variable_to_check_48[1] = enable_variable_46_to_check_48;

// 拆分后校验节点48传递给变量节点87的值以及对变量节点87传递过来的值
wire [5:0] value_check_48_to_variable_87;
wire enable_check_48_to_variable_87;
wire [5:0] value_variable_87_to_check_48;
wire enable_variable_87_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_87 = value_check_48_to_variable[17:12];
assign enable_check_48_to_variable_87 = enable_check_48_to_variable[2];
// 对变量节点87传递过来的值进行组合
assign value_variable_to_check_48[17:12] = value_variable_87_to_check_48;
assign enable_variable_to_check_48[2] = enable_variable_87_to_check_48;

// 拆分后校验节点48传递给变量节点160的值以及对变量节点160传递过来的值
wire [5:0] value_check_48_to_variable_160;
wire enable_check_48_to_variable_160;
wire [5:0] value_variable_160_to_check_48;
wire enable_variable_160_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_160 = value_check_48_to_variable[23:18];
assign enable_check_48_to_variable_160 = enable_check_48_to_variable[3];
// 对变量节点160传递过来的值进行组合
assign value_variable_to_check_48[23:18] = value_variable_160_to_check_48;
assign enable_variable_to_check_48[3] = enable_variable_160_to_check_48;

// 拆分后校验节点48传递给变量节点185的值以及对变量节点185传递过来的值
wire [5:0] value_check_48_to_variable_185;
wire enable_check_48_to_variable_185;
wire [5:0] value_variable_185_to_check_48;
wire enable_variable_185_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_185 = value_check_48_to_variable[29:24];
assign enable_check_48_to_variable_185 = enable_check_48_to_variable[4];
// 对变量节点185传递过来的值进行组合
assign value_variable_to_check_48[29:24] = value_variable_185_to_check_48;
assign enable_variable_to_check_48[4] = enable_variable_185_to_check_48;

// 拆分后校验节点48传递给变量节点243的值以及对变量节点243传递过来的值
wire [5:0] value_check_48_to_variable_243;
wire enable_check_48_to_variable_243;
wire [5:0] value_variable_243_to_check_48;
wire enable_variable_243_to_check_48;
// 对校验节点48的输出值进行拆分
assign value_check_48_to_variable_243 = value_check_48_to_variable[35:30];
assign enable_check_48_to_variable_243 = enable_check_48_to_variable[5];
// 对变量节点243传递过来的值进行组合
assign value_variable_to_check_48[35:30] = value_variable_243_to_check_48;
assign enable_variable_to_check_48[5] = enable_variable_243_to_check_48;


// 校验节点49的接口
wire [35:0] value_variable_to_check_49;
wire [35:0] value_check_49_to_variable;
wire [5:0] enable_variable_to_check_49;
wire [5:0] enable_check_49_to_variable;

// 拆分后校验节点49传递给变量节点32的值以及对变量节点32传递过来的值
wire [5:0] value_check_49_to_variable_32;
wire enable_check_49_to_variable_32;
wire [5:0] value_variable_32_to_check_49;
wire enable_variable_32_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_32 = value_check_49_to_variable[5:0];
assign enable_check_49_to_variable_32 = enable_check_49_to_variable[0];
// 对变量节点32传递过来的值进行组合
assign value_variable_to_check_49[5:0] = value_variable_32_to_check_49;
assign enable_variable_to_check_49[0] = enable_variable_32_to_check_49;

// 拆分后校验节点49传递给变量节点74的值以及对变量节点74传递过来的值
wire [5:0] value_check_49_to_variable_74;
wire enable_check_49_to_variable_74;
wire [5:0] value_variable_74_to_check_49;
wire enable_variable_74_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_74 = value_check_49_to_variable[11:6];
assign enable_check_49_to_variable_74 = enable_check_49_to_variable[1];
// 对变量节点74传递过来的值进行组合
assign value_variable_to_check_49[11:6] = value_variable_74_to_check_49;
assign enable_variable_to_check_49[1] = enable_variable_74_to_check_49;

// 拆分后校验节点49传递给变量节点119的值以及对变量节点119传递过来的值
wire [5:0] value_check_49_to_variable_119;
wire enable_check_49_to_variable_119;
wire [5:0] value_variable_119_to_check_49;
wire enable_variable_119_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_119 = value_check_49_to_variable[17:12];
assign enable_check_49_to_variable_119 = enable_check_49_to_variable[2];
// 对变量节点119传递过来的值进行组合
assign value_variable_to_check_49[17:12] = value_variable_119_to_check_49;
assign enable_variable_to_check_49[2] = enable_variable_119_to_check_49;

// 拆分后校验节点49传递给变量节点136的值以及对变量节点136传递过来的值
wire [5:0] value_check_49_to_variable_136;
wire enable_check_49_to_variable_136;
wire [5:0] value_variable_136_to_check_49;
wire enable_variable_136_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_136 = value_check_49_to_variable[23:18];
assign enable_check_49_to_variable_136 = enable_check_49_to_variable[3];
// 对变量节点136传递过来的值进行组合
assign value_variable_to_check_49[23:18] = value_variable_136_to_check_49;
assign enable_variable_to_check_49[3] = enable_variable_136_to_check_49;

// 拆分后校验节点49传递给变量节点183的值以及对变量节点183传递过来的值
wire [5:0] value_check_49_to_variable_183;
wire enable_check_49_to_variable_183;
wire [5:0] value_variable_183_to_check_49;
wire enable_variable_183_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_183 = value_check_49_to_variable[29:24];
assign enable_check_49_to_variable_183 = enable_check_49_to_variable[4];
// 对变量节点183传递过来的值进行组合
assign value_variable_to_check_49[29:24] = value_variable_183_to_check_49;
assign enable_variable_to_check_49[4] = enable_variable_183_to_check_49;

// 拆分后校验节点49传递给变量节点240的值以及对变量节点240传递过来的值
wire [5:0] value_check_49_to_variable_240;
wire enable_check_49_to_variable_240;
wire [5:0] value_variable_240_to_check_49;
wire enable_variable_240_to_check_49;
// 对校验节点49的输出值进行拆分
assign value_check_49_to_variable_240 = value_check_49_to_variable[35:30];
assign enable_check_49_to_variable_240 = enable_check_49_to_variable[5];
// 对变量节点240传递过来的值进行组合
assign value_variable_to_check_49[35:30] = value_variable_240_to_check_49;
assign enable_variable_to_check_49[5] = enable_variable_240_to_check_49;


// 校验节点50的接口
wire [35:0] value_variable_to_check_50;
wire [35:0] value_check_50_to_variable;
wire [5:0] enable_variable_to_check_50;
wire [5:0] enable_check_50_to_variable;

// 拆分后校验节点50传递给变量节点32的值以及对变量节点32传递过来的值
wire [5:0] value_check_50_to_variable_32;
wire enable_check_50_to_variable_32;
wire [5:0] value_variable_32_to_check_50;
wire enable_variable_32_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_32 = value_check_50_to_variable[5:0];
assign enable_check_50_to_variable_32 = enable_check_50_to_variable[0];
// 对变量节点32传递过来的值进行组合
assign value_variable_to_check_50[5:0] = value_variable_32_to_check_50;
assign enable_variable_to_check_50[0] = enable_variable_32_to_check_50;

// 拆分后校验节点50传递给变量节点43的值以及对变量节点43传递过来的值
wire [5:0] value_check_50_to_variable_43;
wire enable_check_50_to_variable_43;
wire [5:0] value_variable_43_to_check_50;
wire enable_variable_43_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_43 = value_check_50_to_variable[11:6];
assign enable_check_50_to_variable_43 = enable_check_50_to_variable[1];
// 对变量节点43传递过来的值进行组合
assign value_variable_to_check_50[11:6] = value_variable_43_to_check_50;
assign enable_variable_to_check_50[1] = enable_variable_43_to_check_50;

// 拆分后校验节点50传递给变量节点104的值以及对变量节点104传递过来的值
wire [5:0] value_check_50_to_variable_104;
wire enable_check_50_to_variable_104;
wire [5:0] value_variable_104_to_check_50;
wire enable_variable_104_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_104 = value_check_50_to_variable[17:12];
assign enable_check_50_to_variable_104 = enable_check_50_to_variable[2];
// 对变量节点104传递过来的值进行组合
assign value_variable_to_check_50[17:12] = value_variable_104_to_check_50;
assign enable_variable_to_check_50[2] = enable_variable_104_to_check_50;

// 拆分后校验节点50传递给变量节点141的值以及对变量节点141传递过来的值
wire [5:0] value_check_50_to_variable_141;
wire enable_check_50_to_variable_141;
wire [5:0] value_variable_141_to_check_50;
wire enable_variable_141_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_141 = value_check_50_to_variable[23:18];
assign enable_check_50_to_variable_141 = enable_check_50_to_variable[3];
// 对变量节点141传递过来的值进行组合
assign value_variable_to_check_50[23:18] = value_variable_141_to_check_50;
assign enable_variable_to_check_50[3] = enable_variable_141_to_check_50;

// 拆分后校验节点50传递给变量节点167的值以及对变量节点167传递过来的值
wire [5:0] value_check_50_to_variable_167;
wire enable_check_50_to_variable_167;
wire [5:0] value_variable_167_to_check_50;
wire enable_variable_167_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_167 = value_check_50_to_variable[29:24];
assign enable_check_50_to_variable_167 = enable_check_50_to_variable[4];
// 对变量节点167传递过来的值进行组合
assign value_variable_to_check_50[29:24] = value_variable_167_to_check_50;
assign enable_variable_to_check_50[4] = enable_variable_167_to_check_50;

// 拆分后校验节点50传递给变量节点235的值以及对变量节点235传递过来的值
wire [5:0] value_check_50_to_variable_235;
wire enable_check_50_to_variable_235;
wire [5:0] value_variable_235_to_check_50;
wire enable_variable_235_to_check_50;
// 对校验节点50的输出值进行拆分
assign value_check_50_to_variable_235 = value_check_50_to_variable[35:30];
assign enable_check_50_to_variable_235 = enable_check_50_to_variable[5];
// 对变量节点235传递过来的值进行组合
assign value_variable_to_check_50[35:30] = value_variable_235_to_check_50;
assign enable_variable_to_check_50[5] = enable_variable_235_to_check_50;


// 校验节点51的接口
wire [35:0] value_variable_to_check_51;
wire [35:0] value_check_51_to_variable;
wire [5:0] enable_variable_to_check_51;
wire [5:0] enable_check_51_to_variable;

// 拆分后校验节点51传递给变量节点7的值以及对变量节点7传递过来的值
wire [5:0] value_check_51_to_variable_7;
wire enable_check_51_to_variable_7;
wire [5:0] value_variable_7_to_check_51;
wire enable_variable_7_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_7 = value_check_51_to_variable[5:0];
assign enable_check_51_to_variable_7 = enable_check_51_to_variable[0];
// 对变量节点7传递过来的值进行组合
assign value_variable_to_check_51[5:0] = value_variable_7_to_check_51;
assign enable_variable_to_check_51[0] = enable_variable_7_to_check_51;

// 拆分后校验节点51传递给变量节点75的值以及对变量节点75传递过来的值
wire [5:0] value_check_51_to_variable_75;
wire enable_check_51_to_variable_75;
wire [5:0] value_variable_75_to_check_51;
wire enable_variable_75_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_75 = value_check_51_to_variable[11:6];
assign enable_check_51_to_variable_75 = enable_check_51_to_variable[1];
// 对变量节点75传递过来的值进行组合
assign value_variable_to_check_51[11:6] = value_variable_75_to_check_51;
assign enable_variable_to_check_51[1] = enable_variable_75_to_check_51;

// 拆分后校验节点51传递给变量节点119的值以及对变量节点119传递过来的值
wire [5:0] value_check_51_to_variable_119;
wire enable_check_51_to_variable_119;
wire [5:0] value_variable_119_to_check_51;
wire enable_variable_119_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_119 = value_check_51_to_variable[17:12];
assign enable_check_51_to_variable_119 = enable_check_51_to_variable[2];
// 对变量节点119传递过来的值进行组合
assign value_variable_to_check_51[17:12] = value_variable_119_to_check_51;
assign enable_variable_to_check_51[2] = enable_variable_119_to_check_51;

// 拆分后校验节点51传递给变量节点150的值以及对变量节点150传递过来的值
wire [5:0] value_check_51_to_variable_150;
wire enable_check_51_to_variable_150;
wire [5:0] value_variable_150_to_check_51;
wire enable_variable_150_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_150 = value_check_51_to_variable[23:18];
assign enable_check_51_to_variable_150 = enable_check_51_to_variable[3];
// 对变量节点150传递过来的值进行组合
assign value_variable_to_check_51[23:18] = value_variable_150_to_check_51;
assign enable_variable_to_check_51[3] = enable_variable_150_to_check_51;

// 拆分后校验节点51传递给变量节点205的值以及对变量节点205传递过来的值
wire [5:0] value_check_51_to_variable_205;
wire enable_check_51_to_variable_205;
wire [5:0] value_variable_205_to_check_51;
wire enable_variable_205_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_205 = value_check_51_to_variable[29:24];
assign enable_check_51_to_variable_205 = enable_check_51_to_variable[4];
// 对变量节点205传递过来的值进行组合
assign value_variable_to_check_51[29:24] = value_variable_205_to_check_51;
assign enable_variable_to_check_51[4] = enable_variable_205_to_check_51;

// 拆分后校验节点51传递给变量节点244的值以及对变量节点244传递过来的值
wire [5:0] value_check_51_to_variable_244;
wire enable_check_51_to_variable_244;
wire [5:0] value_variable_244_to_check_51;
wire enable_variable_244_to_check_51;
// 对校验节点51的输出值进行拆分
assign value_check_51_to_variable_244 = value_check_51_to_variable[35:30];
assign enable_check_51_to_variable_244 = enable_check_51_to_variable[5];
// 对变量节点244传递过来的值进行组合
assign value_variable_to_check_51[35:30] = value_variable_244_to_check_51;
assign enable_variable_to_check_51[5] = enable_variable_244_to_check_51;


// 校验节点52的接口
wire [35:0] value_variable_to_check_52;
wire [35:0] value_check_52_to_variable;
wire [5:0] enable_variable_to_check_52;
wire [5:0] enable_check_52_to_variable;

// 拆分后校验节点52传递给变量节点32的值以及对变量节点32传递过来的值
wire [5:0] value_check_52_to_variable_32;
wire enable_check_52_to_variable_32;
wire [5:0] value_variable_32_to_check_52;
wire enable_variable_32_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_32 = value_check_52_to_variable[5:0];
assign enable_check_52_to_variable_32 = enable_check_52_to_variable[0];
// 对变量节点32传递过来的值进行组合
assign value_variable_to_check_52[5:0] = value_variable_32_to_check_52;
assign enable_variable_to_check_52[0] = enable_variable_32_to_check_52;

// 拆分后校验节点52传递给变量节点58的值以及对变量节点58传递过来的值
wire [5:0] value_check_52_to_variable_58;
wire enable_check_52_to_variable_58;
wire [5:0] value_variable_58_to_check_52;
wire enable_variable_58_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_58 = value_check_52_to_variable[11:6];
assign enable_check_52_to_variable_58 = enable_check_52_to_variable[1];
// 对变量节点58传递过来的值进行组合
assign value_variable_to_check_52[11:6] = value_variable_58_to_check_52;
assign enable_variable_to_check_52[1] = enable_variable_58_to_check_52;

// 拆分后校验节点52传递给变量节点120的值以及对变量节点120传递过来的值
wire [5:0] value_check_52_to_variable_120;
wire enable_check_52_to_variable_120;
wire [5:0] value_variable_120_to_check_52;
wire enable_variable_120_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_120 = value_check_52_to_variable[17:12];
assign enable_check_52_to_variable_120 = enable_check_52_to_variable[2];
// 对变量节点120传递过来的值进行组合
assign value_variable_to_check_52[17:12] = value_variable_120_to_check_52;
assign enable_variable_to_check_52[2] = enable_variable_120_to_check_52;

// 拆分后校验节点52传递给变量节点161的值以及对变量节点161传递过来的值
wire [5:0] value_check_52_to_variable_161;
wire enable_check_52_to_variable_161;
wire [5:0] value_variable_161_to_check_52;
wire enable_variable_161_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_161 = value_check_52_to_variable[23:18];
assign enable_check_52_to_variable_161 = enable_check_52_to_variable[3];
// 对变量节点161传递过来的值进行组合
assign value_variable_to_check_52[23:18] = value_variable_161_to_check_52;
assign enable_variable_to_check_52[3] = enable_variable_161_to_check_52;

// 拆分后校验节点52传递给变量节点182的值以及对变量节点182传递过来的值
wire [5:0] value_check_52_to_variable_182;
wire enable_check_52_to_variable_182;
wire [5:0] value_variable_182_to_check_52;
wire enable_variable_182_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_182 = value_check_52_to_variable[29:24];
assign enable_check_52_to_variable_182 = enable_check_52_to_variable[4];
// 对变量节点182传递过来的值进行组合
assign value_variable_to_check_52[29:24] = value_variable_182_to_check_52;
assign enable_variable_to_check_52[4] = enable_variable_182_to_check_52;

// 拆分后校验节点52传递给变量节点231的值以及对变量节点231传递过来的值
wire [5:0] value_check_52_to_variable_231;
wire enable_check_52_to_variable_231;
wire [5:0] value_variable_231_to_check_52;
wire enable_variable_231_to_check_52;
// 对校验节点52的输出值进行拆分
assign value_check_52_to_variable_231 = value_check_52_to_variable[35:30];
assign enable_check_52_to_variable_231 = enable_check_52_to_variable[5];
// 对变量节点231传递过来的值进行组合
assign value_variable_to_check_52[35:30] = value_variable_231_to_check_52;
assign enable_variable_to_check_52[5] = enable_variable_231_to_check_52;


// 校验节点53的接口
wire [35:0] value_variable_to_check_53;
wire [35:0] value_check_53_to_variable;
wire [5:0] enable_variable_to_check_53;
wire [5:0] enable_check_53_to_variable;

// 拆分后校验节点53传递给变量节点33的值以及对变量节点33传递过来的值
wire [5:0] value_check_53_to_variable_33;
wire enable_check_53_to_variable_33;
wire [5:0] value_variable_33_to_check_53;
wire enable_variable_33_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_33 = value_check_53_to_variable[5:0];
assign enable_check_53_to_variable_33 = enable_check_53_to_variable[0];
// 对变量节点33传递过来的值进行组合
assign value_variable_to_check_53[5:0] = value_variable_33_to_check_53;
assign enable_variable_to_check_53[0] = enable_variable_33_to_check_53;

// 拆分后校验节点53传递给变量节点63的值以及对变量节点63传递过来的值
wire [5:0] value_check_53_to_variable_63;
wire enable_check_53_to_variable_63;
wire [5:0] value_variable_63_to_check_53;
wire enable_variable_63_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_63 = value_check_53_to_variable[11:6];
assign enable_check_53_to_variable_63 = enable_check_53_to_variable[1];
// 对变量节点63传递过来的值进行组合
assign value_variable_to_check_53[11:6] = value_variable_63_to_check_53;
assign enable_variable_to_check_53[1] = enable_variable_63_to_check_53;

// 拆分后校验节点53传递给变量节点121的值以及对变量节点121传递过来的值
wire [5:0] value_check_53_to_variable_121;
wire enable_check_53_to_variable_121;
wire [5:0] value_variable_121_to_check_53;
wire enable_variable_121_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_121 = value_check_53_to_variable[17:12];
assign enable_check_53_to_variable_121 = enable_check_53_to_variable[2];
// 对变量节点121传递过来的值进行组合
assign value_variable_to_check_53[17:12] = value_variable_121_to_check_53;
assign enable_variable_to_check_53[2] = enable_variable_121_to_check_53;

// 拆分后校验节点53传递给变量节点152的值以及对变量节点152传递过来的值
wire [5:0] value_check_53_to_variable_152;
wire enable_check_53_to_variable_152;
wire [5:0] value_variable_152_to_check_53;
wire enable_variable_152_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_152 = value_check_53_to_variable[23:18];
assign enable_check_53_to_variable_152 = enable_check_53_to_variable[3];
// 对变量节点152传递过来的值进行组合
assign value_variable_to_check_53[23:18] = value_variable_152_to_check_53;
assign enable_variable_to_check_53[3] = enable_variable_152_to_check_53;

// 拆分后校验节点53传递给变量节点174的值以及对变量节点174传递过来的值
wire [5:0] value_check_53_to_variable_174;
wire enable_check_53_to_variable_174;
wire [5:0] value_variable_174_to_check_53;
wire enable_variable_174_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_174 = value_check_53_to_variable[29:24];
assign enable_check_53_to_variable_174 = enable_check_53_to_variable[4];
// 对变量节点174传递过来的值进行组合
assign value_variable_to_check_53[29:24] = value_variable_174_to_check_53;
assign enable_variable_to_check_53[4] = enable_variable_174_to_check_53;

// 拆分后校验节点53传递给变量节点243的值以及对变量节点243传递过来的值
wire [5:0] value_check_53_to_variable_243;
wire enable_check_53_to_variable_243;
wire [5:0] value_variable_243_to_check_53;
wire enable_variable_243_to_check_53;
// 对校验节点53的输出值进行拆分
assign value_check_53_to_variable_243 = value_check_53_to_variable[35:30];
assign enable_check_53_to_variable_243 = enable_check_53_to_variable[5];
// 对变量节点243传递过来的值进行组合
assign value_variable_to_check_53[35:30] = value_variable_243_to_check_53;
assign enable_variable_to_check_53[5] = enable_variable_243_to_check_53;


// 校验节点54的接口
wire [35:0] value_variable_to_check_54;
wire [35:0] value_check_54_to_variable;
wire [5:0] enable_variable_to_check_54;
wire [5:0] enable_check_54_to_variable;

// 拆分后校验节点54传递给变量节点31的值以及对变量节点31传递过来的值
wire [5:0] value_check_54_to_variable_31;
wire enable_check_54_to_variable_31;
wire [5:0] value_variable_31_to_check_54;
wire enable_variable_31_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_31 = value_check_54_to_variable[5:0];
assign enable_check_54_to_variable_31 = enable_check_54_to_variable[0];
// 对变量节点31传递过来的值进行组合
assign value_variable_to_check_54[5:0] = value_variable_31_to_check_54;
assign enable_variable_to_check_54[0] = enable_variable_31_to_check_54;

// 拆分后校验节点54传递给变量节点45的值以及对变量节点45传递过来的值
wire [5:0] value_check_54_to_variable_45;
wire enable_check_54_to_variable_45;
wire [5:0] value_variable_45_to_check_54;
wire enable_variable_45_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_45 = value_check_54_to_variable[11:6];
assign enable_check_54_to_variable_45 = enable_check_54_to_variable[1];
// 对变量节点45传递过来的值进行组合
assign value_variable_to_check_54[11:6] = value_variable_45_to_check_54;
assign enable_variable_to_check_54[1] = enable_variable_45_to_check_54;

// 拆分后校验节点54传递给变量节点106的值以及对变量节点106传递过来的值
wire [5:0] value_check_54_to_variable_106;
wire enable_check_54_to_variable_106;
wire [5:0] value_variable_106_to_check_54;
wire enable_variable_106_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_106 = value_check_54_to_variable[17:12];
assign enable_check_54_to_variable_106 = enable_check_54_to_variable[2];
// 对变量节点106传递过来的值进行组合
assign value_variable_to_check_54[17:12] = value_variable_106_to_check_54;
assign enable_variable_to_check_54[2] = enable_variable_106_to_check_54;

// 拆分后校验节点54传递给变量节点162的值以及对变量节点162传递过来的值
wire [5:0] value_check_54_to_variable_162;
wire enable_check_54_to_variable_162;
wire [5:0] value_variable_162_to_check_54;
wire enable_variable_162_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_162 = value_check_54_to_variable[23:18];
assign enable_check_54_to_variable_162 = enable_check_54_to_variable[3];
// 对变量节点162传递过来的值进行组合
assign value_variable_to_check_54[23:18] = value_variable_162_to_check_54;
assign enable_variable_to_check_54[3] = enable_variable_162_to_check_54;

// 拆分后校验节点54传递给变量节点193的值以及对变量节点193传递过来的值
wire [5:0] value_check_54_to_variable_193;
wire enable_check_54_to_variable_193;
wire [5:0] value_variable_193_to_check_54;
wire enable_variable_193_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_193 = value_check_54_to_variable[29:24];
assign enable_check_54_to_variable_193 = enable_check_54_to_variable[4];
// 对变量节点193传递过来的值进行组合
assign value_variable_to_check_54[29:24] = value_variable_193_to_check_54;
assign enable_variable_to_check_54[4] = enable_variable_193_to_check_54;

// 拆分后校验节点54传递给变量节点233的值以及对变量节点233传递过来的值
wire [5:0] value_check_54_to_variable_233;
wire enable_check_54_to_variable_233;
wire [5:0] value_variable_233_to_check_54;
wire enable_variable_233_to_check_54;
// 对校验节点54的输出值进行拆分
assign value_check_54_to_variable_233 = value_check_54_to_variable[35:30];
assign enable_check_54_to_variable_233 = enable_check_54_to_variable[5];
// 对变量节点233传递过来的值进行组合
assign value_variable_to_check_54[35:30] = value_variable_233_to_check_54;
assign enable_variable_to_check_54[5] = enable_variable_233_to_check_54;


// 校验节点55的接口
wire [35:0] value_variable_to_check_55;
wire [35:0] value_check_55_to_variable;
wire [5:0] enable_variable_to_check_55;
wire [5:0] enable_check_55_to_variable;

// 拆分后校验节点55传递给变量节点34的值以及对变量节点34传递过来的值
wire [5:0] value_check_55_to_variable_34;
wire enable_check_55_to_variable_34;
wire [5:0] value_variable_34_to_check_55;
wire enable_variable_34_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_34 = value_check_55_to_variable[5:0];
assign enable_check_55_to_variable_34 = enable_check_55_to_variable[0];
// 对变量节点34传递过来的值进行组合
assign value_variable_to_check_55[5:0] = value_variable_34_to_check_55;
assign enable_variable_to_check_55[0] = enable_variable_34_to_check_55;

// 拆分后校验节点55传递给变量节点62的值以及对变量节点62传递过来的值
wire [5:0] value_check_55_to_variable_62;
wire enable_check_55_to_variable_62;
wire [5:0] value_variable_62_to_check_55;
wire enable_variable_62_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_62 = value_check_55_to_variable[11:6];
assign enable_check_55_to_variable_62 = enable_check_55_to_variable[1];
// 对变量节点62传递过来的值进行组合
assign value_variable_to_check_55[11:6] = value_variable_62_to_check_55;
assign enable_variable_to_check_55[1] = enable_variable_62_to_check_55;

// 拆分后校验节点55传递给变量节点103的值以及对变量节点103传递过来的值
wire [5:0] value_check_55_to_variable_103;
wire enable_check_55_to_variable_103;
wire [5:0] value_variable_103_to_check_55;
wire enable_variable_103_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_103 = value_check_55_to_variable[17:12];
assign enable_check_55_to_variable_103 = enable_check_55_to_variable[2];
// 对变量节点103传递过来的值进行组合
assign value_variable_to_check_55[17:12] = value_variable_103_to_check_55;
assign enable_variable_to_check_55[2] = enable_variable_103_to_check_55;

// 拆分后校验节点55传递给变量节点134的值以及对变量节点134传递过来的值
wire [5:0] value_check_55_to_variable_134;
wire enable_check_55_to_variable_134;
wire [5:0] value_variable_134_to_check_55;
wire enable_variable_134_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_134 = value_check_55_to_variable[23:18];
assign enable_check_55_to_variable_134 = enable_check_55_to_variable[3];
// 对变量节点134传递过来的值进行组合
assign value_variable_to_check_55[23:18] = value_variable_134_to_check_55;
assign enable_variable_to_check_55[3] = enable_variable_134_to_check_55;

// 拆分后校验节点55传递给变量节点177的值以及对变量节点177传递过来的值
wire [5:0] value_check_55_to_variable_177;
wire enable_check_55_to_variable_177;
wire [5:0] value_variable_177_to_check_55;
wire enable_variable_177_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_177 = value_check_55_to_variable[29:24];
assign enable_check_55_to_variable_177 = enable_check_55_to_variable[4];
// 对变量节点177传递过来的值进行组合
assign value_variable_to_check_55[29:24] = value_variable_177_to_check_55;
assign enable_variable_to_check_55[4] = enable_variable_177_to_check_55;

// 拆分后校验节点55传递给变量节点245的值以及对变量节点245传递过来的值
wire [5:0] value_check_55_to_variable_245;
wire enable_check_55_to_variable_245;
wire [5:0] value_variable_245_to_check_55;
wire enable_variable_245_to_check_55;
// 对校验节点55的输出值进行拆分
assign value_check_55_to_variable_245 = value_check_55_to_variable[35:30];
assign enable_check_55_to_variable_245 = enable_check_55_to_variable[5];
// 对变量节点245传递过来的值进行组合
assign value_variable_to_check_55[35:30] = value_variable_245_to_check_55;
assign enable_variable_to_check_55[5] = enable_variable_245_to_check_55;


// 校验节点56的接口
wire [35:0] value_variable_to_check_56;
wire [35:0] value_check_56_to_variable;
wire [5:0] enable_variable_to_check_56;
wire [5:0] enable_check_56_to_variable;

// 拆分后校验节点56传递给变量节点18的值以及对变量节点18传递过来的值
wire [5:0] value_check_56_to_variable_18;
wire enable_check_56_to_variable_18;
wire [5:0] value_variable_18_to_check_56;
wire enable_variable_18_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_18 = value_check_56_to_variable[5:0];
assign enable_check_56_to_variable_18 = enable_check_56_to_variable[0];
// 对变量节点18传递过来的值进行组合
assign value_variable_to_check_56[5:0] = value_variable_18_to_check_56;
assign enable_variable_to_check_56[0] = enable_variable_18_to_check_56;

// 拆分后校验节点56传递给变量节点60的值以及对变量节点60传递过来的值
wire [5:0] value_check_56_to_variable_60;
wire enable_check_56_to_variable_60;
wire [5:0] value_variable_60_to_check_56;
wire enable_variable_60_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_60 = value_check_56_to_variable[11:6];
assign enable_check_56_to_variable_60 = enable_check_56_to_variable[1];
// 对变量节点60传递过来的值进行组合
assign value_variable_to_check_56[11:6] = value_variable_60_to_check_56;
assign enable_variable_to_check_56[1] = enable_variable_60_to_check_56;

// 拆分后校验节点56传递给变量节点117的值以及对变量节点117传递过来的值
wire [5:0] value_check_56_to_variable_117;
wire enable_check_56_to_variable_117;
wire [5:0] value_variable_117_to_check_56;
wire enable_variable_117_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_117 = value_check_56_to_variable[17:12];
assign enable_check_56_to_variable_117 = enable_check_56_to_variable[2];
// 对变量节点117传递过来的值进行组合
assign value_variable_to_check_56[17:12] = value_variable_117_to_check_56;
assign enable_variable_to_check_56[2] = enable_variable_117_to_check_56;

// 拆分后校验节点56传递给变量节点163的值以及对变量节点163传递过来的值
wire [5:0] value_check_56_to_variable_163;
wire enable_check_56_to_variable_163;
wire [5:0] value_variable_163_to_check_56;
wire enable_variable_163_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_163 = value_check_56_to_variable[23:18];
assign enable_check_56_to_variable_163 = enable_check_56_to_variable[3];
// 对变量节点163传递过来的值进行组合
assign value_variable_to_check_56[23:18] = value_variable_163_to_check_56;
assign enable_variable_to_check_56[3] = enable_variable_163_to_check_56;

// 拆分后校验节点56传递给变量节点206的值以及对变量节点206传递过来的值
wire [5:0] value_check_56_to_variable_206;
wire enable_check_56_to_variable_206;
wire [5:0] value_variable_206_to_check_56;
wire enable_variable_206_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_206 = value_check_56_to_variable[29:24];
assign enable_check_56_to_variable_206 = enable_check_56_to_variable[4];
// 对变量节点206传递过来的值进行组合
assign value_variable_to_check_56[29:24] = value_variable_206_to_check_56;
assign enable_variable_to_check_56[4] = enable_variable_206_to_check_56;

// 拆分后校验节点56传递给变量节点224的值以及对变量节点224传递过来的值
wire [5:0] value_check_56_to_variable_224;
wire enable_check_56_to_variable_224;
wire [5:0] value_variable_224_to_check_56;
wire enable_variable_224_to_check_56;
// 对校验节点56的输出值进行拆分
assign value_check_56_to_variable_224 = value_check_56_to_variable[35:30];
assign enable_check_56_to_variable_224 = enable_check_56_to_variable[5];
// 对变量节点224传递过来的值进行组合
assign value_variable_to_check_56[35:30] = value_variable_224_to_check_56;
assign enable_variable_to_check_56[5] = enable_variable_224_to_check_56;


// 校验节点57的接口
wire [35:0] value_variable_to_check_57;
wire [35:0] value_check_57_to_variable;
wire [5:0] enable_variable_to_check_57;
wire [5:0] enable_check_57_to_variable;

// 拆分后校验节点57传递给变量节点8的值以及对变量节点8传递过来的值
wire [5:0] value_check_57_to_variable_8;
wire enable_check_57_to_variable_8;
wire [5:0] value_variable_8_to_check_57;
wire enable_variable_8_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_8 = value_check_57_to_variable[5:0];
assign enable_check_57_to_variable_8 = enable_check_57_to_variable[0];
// 对变量节点8传递过来的值进行组合
assign value_variable_to_check_57[5:0] = value_variable_8_to_check_57;
assign enable_variable_to_check_57[0] = enable_variable_8_to_check_57;

// 拆分后校验节点57传递给变量节点76的值以及对变量节点76传递过来的值
wire [5:0] value_check_57_to_variable_76;
wire enable_check_57_to_variable_76;
wire [5:0] value_variable_76_to_check_57;
wire enable_variable_76_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_76 = value_check_57_to_variable[11:6];
assign enable_check_57_to_variable_76 = enable_check_57_to_variable[1];
// 对变量节点76传递过来的值进行组合
assign value_variable_to_check_57[11:6] = value_variable_76_to_check_57;
assign enable_variable_to_check_57[1] = enable_variable_76_to_check_57;

// 拆分后校验节点57传递给变量节点86的值以及对变量节点86传递过来的值
wire [5:0] value_check_57_to_variable_86;
wire enable_check_57_to_variable_86;
wire [5:0] value_variable_86_to_check_57;
wire enable_variable_86_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_86 = value_check_57_to_variable[17:12];
assign enable_check_57_to_variable_86 = enable_check_57_to_variable[2];
// 对变量节点86传递过来的值进行组合
assign value_variable_to_check_57[17:12] = value_variable_86_to_check_57;
assign enable_variable_to_check_57[2] = enable_variable_86_to_check_57;

// 拆分后校验节点57传递给变量节点100的值以及对变量节点100传递过来的值
wire [5:0] value_check_57_to_variable_100;
wire enable_check_57_to_variable_100;
wire [5:0] value_variable_100_to_check_57;
wire enable_variable_100_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_100 = value_check_57_to_variable[23:18];
assign enable_check_57_to_variable_100 = enable_check_57_to_variable[3];
// 对变量节点100传递过来的值进行组合
assign value_variable_to_check_57[23:18] = value_variable_100_to_check_57;
assign enable_variable_to_check_57[3] = enable_variable_100_to_check_57;

// 拆分后校验节点57传递给变量节点172的值以及对变量节点172传递过来的值
wire [5:0] value_check_57_to_variable_172;
wire enable_check_57_to_variable_172;
wire [5:0] value_variable_172_to_check_57;
wire enable_variable_172_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_172 = value_check_57_to_variable[29:24];
assign enable_check_57_to_variable_172 = enable_check_57_to_variable[4];
// 对变量节点172传递过来的值进行组合
assign value_variable_to_check_57[29:24] = value_variable_172_to_check_57;
assign enable_variable_to_check_57[4] = enable_variable_172_to_check_57;

// 拆分后校验节点57传递给变量节点228的值以及对变量节点228传递过来的值
wire [5:0] value_check_57_to_variable_228;
wire enable_check_57_to_variable_228;
wire [5:0] value_variable_228_to_check_57;
wire enable_variable_228_to_check_57;
// 对校验节点57的输出值进行拆分
assign value_check_57_to_variable_228 = value_check_57_to_variable[35:30];
assign enable_check_57_to_variable_228 = enable_check_57_to_variable[5];
// 对变量节点228传递过来的值进行组合
assign value_variable_to_check_57[35:30] = value_variable_228_to_check_57;
assign enable_variable_to_check_57[5] = enable_variable_228_to_check_57;


// 校验节点58的接口
wire [35:0] value_variable_to_check_58;
wire [35:0] value_check_58_to_variable;
wire [5:0] enable_variable_to_check_58;
wire [5:0] enable_check_58_to_variable;

// 拆分后校验节点58传递给变量节点35的值以及对变量节点35传递过来的值
wire [5:0] value_check_58_to_variable_35;
wire enable_check_58_to_variable_35;
wire [5:0] value_variable_35_to_check_58;
wire enable_variable_35_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_35 = value_check_58_to_variable[5:0];
assign enable_check_58_to_variable_35 = enable_check_58_to_variable[0];
// 对变量节点35传递过来的值进行组合
assign value_variable_to_check_58[5:0] = value_variable_35_to_check_58;
assign enable_variable_to_check_58[0] = enable_variable_35_to_check_58;

// 拆分后校验节点58传递给变量节点73的值以及对变量节点73传递过来的值
wire [5:0] value_check_58_to_variable_73;
wire enable_check_58_to_variable_73;
wire [5:0] value_variable_73_to_check_58;
wire enable_variable_73_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_73 = value_check_58_to_variable[11:6];
assign enable_check_58_to_variable_73 = enable_check_58_to_variable[1];
// 对变量节点73传递过来的值进行组合
assign value_variable_to_check_58[11:6] = value_variable_73_to_check_58;
assign enable_variable_to_check_58[1] = enable_variable_73_to_check_58;

// 拆分后校验节点58传递给变量节点109的值以及对变量节点109传递过来的值
wire [5:0] value_check_58_to_variable_109;
wire enable_check_58_to_variable_109;
wire [5:0] value_variable_109_to_check_58;
wire enable_variable_109_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_109 = value_check_58_to_variable[17:12];
assign enable_check_58_to_variable_109 = enable_check_58_to_variable[2];
// 对变量节点109传递过来的值进行组合
assign value_variable_to_check_58[17:12] = value_variable_109_to_check_58;
assign enable_variable_to_check_58[2] = enable_variable_109_to_check_58;

// 拆分后校验节点58传递给变量节点138的值以及对变量节点138传递过来的值
wire [5:0] value_check_58_to_variable_138;
wire enable_check_58_to_variable_138;
wire [5:0] value_variable_138_to_check_58;
wire enable_variable_138_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_138 = value_check_58_to_variable[23:18];
assign enable_check_58_to_variable_138 = enable_check_58_to_variable[3];
// 对变量节点138传递过来的值进行组合
assign value_variable_to_check_58[23:18] = value_variable_138_to_check_58;
assign enable_variable_to_check_58[3] = enable_variable_138_to_check_58;

// 拆分后校验节点58传递给变量节点204的值以及对变量节点204传递过来的值
wire [5:0] value_check_58_to_variable_204;
wire enable_check_58_to_variable_204;
wire [5:0] value_variable_204_to_check_58;
wire enable_variable_204_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_204 = value_check_58_to_variable[29:24];
assign enable_check_58_to_variable_204 = enable_check_58_to_variable[4];
// 对变量节点204传递过来的值进行组合
assign value_variable_to_check_58[29:24] = value_variable_204_to_check_58;
assign enable_variable_to_check_58[4] = enable_variable_204_to_check_58;

// 拆分后校验节点58传递给变量节点246的值以及对变量节点246传递过来的值
wire [5:0] value_check_58_to_variable_246;
wire enable_check_58_to_variable_246;
wire [5:0] value_variable_246_to_check_58;
wire enable_variable_246_to_check_58;
// 对校验节点58的输出值进行拆分
assign value_check_58_to_variable_246 = value_check_58_to_variable[35:30];
assign enable_check_58_to_variable_246 = enable_check_58_to_variable[5];
// 对变量节点246传递过来的值进行组合
assign value_variable_to_check_58[35:30] = value_variable_246_to_check_58;
assign enable_variable_to_check_58[5] = enable_variable_246_to_check_58;


// 校验节点59的接口
wire [35:0] value_variable_to_check_59;
wire [35:0] value_check_59_to_variable;
wire [5:0] enable_variable_to_check_59;
wire [5:0] enable_check_59_to_variable;

// 拆分后校验节点59传递给变量节点24的值以及对变量节点24传递过来的值
wire [5:0] value_check_59_to_variable_24;
wire enable_check_59_to_variable_24;
wire [5:0] value_variable_24_to_check_59;
wire enable_variable_24_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_24 = value_check_59_to_variable[5:0];
assign enable_check_59_to_variable_24 = enable_check_59_to_variable[0];
// 对变量节点24传递过来的值进行组合
assign value_variable_to_check_59[5:0] = value_variable_24_to_check_59;
assign enable_variable_to_check_59[0] = enable_variable_24_to_check_59;

// 拆分后校验节点59传递给变量节点77的值以及对变量节点77传递过来的值
wire [5:0] value_check_59_to_variable_77;
wire enable_check_59_to_variable_77;
wire [5:0] value_variable_77_to_check_59;
wire enable_variable_77_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_77 = value_check_59_to_variable[11:6];
assign enable_check_59_to_variable_77 = enable_check_59_to_variable[1];
// 对变量节点77传递过来的值进行组合
assign value_variable_to_check_59[11:6] = value_variable_77_to_check_59;
assign enable_variable_to_check_59[1] = enable_variable_77_to_check_59;

// 拆分后校验节点59传递给变量节点99的值以及对变量节点99传递过来的值
wire [5:0] value_check_59_to_variable_99;
wire enable_check_59_to_variable_99;
wire [5:0] value_variable_99_to_check_59;
wire enable_variable_99_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_99 = value_check_59_to_variable[17:12];
assign enable_check_59_to_variable_99 = enable_check_59_to_variable[2];
// 对变量节点99传递过来的值进行组合
assign value_variable_to_check_59[17:12] = value_variable_99_to_check_59;
assign enable_variable_to_check_59[2] = enable_variable_99_to_check_59;

// 拆分后校验节点59传递给变量节点146的值以及对变量节点146传递过来的值
wire [5:0] value_check_59_to_variable_146;
wire enable_check_59_to_variable_146;
wire [5:0] value_variable_146_to_check_59;
wire enable_variable_146_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_146 = value_check_59_to_variable[23:18];
assign enable_check_59_to_variable_146 = enable_check_59_to_variable[3];
// 对变量节点146传递过来的值进行组合
assign value_variable_to_check_59[23:18] = value_variable_146_to_check_59;
assign enable_variable_to_check_59[3] = enable_variable_146_to_check_59;

// 拆分后校验节点59传递给变量节点193的值以及对变量节点193传递过来的值
wire [5:0] value_check_59_to_variable_193;
wire enable_check_59_to_variable_193;
wire [5:0] value_variable_193_to_check_59;
wire enable_variable_193_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_193 = value_check_59_to_variable[29:24];
assign enable_check_59_to_variable_193 = enable_check_59_to_variable[4];
// 对变量节点193传递过来的值进行组合
assign value_variable_to_check_59[29:24] = value_variable_193_to_check_59;
assign enable_variable_to_check_59[4] = enable_variable_193_to_check_59;

// 拆分后校验节点59传递给变量节点246的值以及对变量节点246传递过来的值
wire [5:0] value_check_59_to_variable_246;
wire enable_check_59_to_variable_246;
wire [5:0] value_variable_246_to_check_59;
wire enable_variable_246_to_check_59;
// 对校验节点59的输出值进行拆分
assign value_check_59_to_variable_246 = value_check_59_to_variable[35:30];
assign enable_check_59_to_variable_246 = enable_check_59_to_variable[5];
// 对变量节点246传递过来的值进行组合
assign value_variable_to_check_59[35:30] = value_variable_246_to_check_59;
assign enable_variable_to_check_59[5] = enable_variable_246_to_check_59;


// 校验节点60的接口
wire [35:0] value_variable_to_check_60;
wire [35:0] value_check_60_to_variable;
wire [5:0] enable_variable_to_check_60;
wire [5:0] enable_check_60_to_variable;

// 拆分后校验节点60传递给变量节点36的值以及对变量节点36传递过来的值
wire [5:0] value_check_60_to_variable_36;
wire enable_check_60_to_variable_36;
wire [5:0] value_variable_36_to_check_60;
wire enable_variable_36_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_36 = value_check_60_to_variable[5:0];
assign enable_check_60_to_variable_36 = enable_check_60_to_variable[0];
// 对变量节点36传递过来的值进行组合
assign value_variable_to_check_60[5:0] = value_variable_36_to_check_60;
assign enable_variable_to_check_60[0] = enable_variable_36_to_check_60;

// 拆分后校验节点60传递给变量节点60的值以及对变量节点60传递过来的值
wire [5:0] value_check_60_to_variable_60;
wire enable_check_60_to_variable_60;
wire [5:0] value_variable_60_to_check_60;
wire enable_variable_60_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_60 = value_check_60_to_variable[11:6];
assign enable_check_60_to_variable_60 = enable_check_60_to_variable[1];
// 对变量节点60传递过来的值进行组合
assign value_variable_to_check_60[11:6] = value_variable_60_to_check_60;
assign enable_variable_to_check_60[1] = enable_variable_60_to_check_60;

// 拆分后校验节点60传递给变量节点122的值以及对变量节点122传递过来的值
wire [5:0] value_check_60_to_variable_122;
wire enable_check_60_to_variable_122;
wire [5:0] value_variable_122_to_check_60;
wire enable_variable_122_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_122 = value_check_60_to_variable[17:12];
assign enable_check_60_to_variable_122 = enable_check_60_to_variable[2];
// 对变量节点122传递过来的值进行组合
assign value_variable_to_check_60[17:12] = value_variable_122_to_check_60;
assign enable_variable_to_check_60[2] = enable_variable_122_to_check_60;

// 拆分后校验节点60传递给变量节点149的值以及对变量节点149传递过来的值
wire [5:0] value_check_60_to_variable_149;
wire enable_check_60_to_variable_149;
wire [5:0] value_variable_149_to_check_60;
wire enable_variable_149_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_149 = value_check_60_to_variable[23:18];
assign enable_check_60_to_variable_149 = enable_check_60_to_variable[3];
// 对变量节点149传递过来的值进行组合
assign value_variable_to_check_60[23:18] = value_variable_149_to_check_60;
assign enable_variable_to_check_60[3] = enable_variable_149_to_check_60;

// 拆分后校验节点60传递给变量节点173的值以及对变量节点173传递过来的值
wire [5:0] value_check_60_to_variable_173;
wire enable_check_60_to_variable_173;
wire [5:0] value_variable_173_to_check_60;
wire enable_variable_173_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_173 = value_check_60_to_variable[29:24];
assign enable_check_60_to_variable_173 = enable_check_60_to_variable[4];
// 对变量节点173传递过来的值进行组合
assign value_variable_to_check_60[29:24] = value_variable_173_to_check_60;
assign enable_variable_to_check_60[4] = enable_variable_173_to_check_60;

// 拆分后校验节点60传递给变量节点247的值以及对变量节点247传递过来的值
wire [5:0] value_check_60_to_variable_247;
wire enable_check_60_to_variable_247;
wire [5:0] value_variable_247_to_check_60;
wire enable_variable_247_to_check_60;
// 对校验节点60的输出值进行拆分
assign value_check_60_to_variable_247 = value_check_60_to_variable[35:30];
assign enable_check_60_to_variable_247 = enable_check_60_to_variable[5];
// 对变量节点247传递过来的值进行组合
assign value_variable_to_check_60[35:30] = value_variable_247_to_check_60;
assign enable_variable_to_check_60[5] = enable_variable_247_to_check_60;


// 校验节点61的接口
wire [35:0] value_variable_to_check_61;
wire [35:0] value_check_61_to_variable;
wire [5:0] enable_variable_to_check_61;
wire [5:0] enable_check_61_to_variable;

// 拆分后校验节点61传递给变量节点7的值以及对变量节点7传递过来的值
wire [5:0] value_check_61_to_variable_7;
wire enable_check_61_to_variable_7;
wire [5:0] value_variable_7_to_check_61;
wire enable_variable_7_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_7 = value_check_61_to_variable[5:0];
assign enable_check_61_to_variable_7 = enable_check_61_to_variable[0];
// 对变量节点7传递过来的值进行组合
assign value_variable_to_check_61[5:0] = value_variable_7_to_check_61;
assign enable_variable_to_check_61[0] = enable_variable_7_to_check_61;

// 拆分后校验节点61传递给变量节点44的值以及对变量节点44传递过来的值
wire [5:0] value_check_61_to_variable_44;
wire enable_check_61_to_variable_44;
wire [5:0] value_variable_44_to_check_61;
wire enable_variable_44_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_44 = value_check_61_to_variable[11:6];
assign enable_check_61_to_variable_44 = enable_check_61_to_variable[1];
// 对变量节点44传递过来的值进行组合
assign value_variable_to_check_61[11:6] = value_variable_44_to_check_61;
assign enable_variable_to_check_61[1] = enable_variable_44_to_check_61;

// 拆分后校验节点61传递给变量节点114的值以及对变量节点114传递过来的值
wire [5:0] value_check_61_to_variable_114;
wire enable_check_61_to_variable_114;
wire [5:0] value_variable_114_to_check_61;
wire enable_variable_114_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_114 = value_check_61_to_variable[17:12];
assign enable_check_61_to_variable_114 = enable_check_61_to_variable[2];
// 对变量节点114传递过来的值进行组合
assign value_variable_to_check_61[17:12] = value_variable_114_to_check_61;
assign enable_variable_to_check_61[2] = enable_variable_114_to_check_61;

// 拆分后校验节点61传递给变量节点151的值以及对变量节点151传递过来的值
wire [5:0] value_check_61_to_variable_151;
wire enable_check_61_to_variable_151;
wire [5:0] value_variable_151_to_check_61;
wire enable_variable_151_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_151 = value_check_61_to_variable[23:18];
assign enable_check_61_to_variable_151 = enable_check_61_to_variable[3];
// 对变量节点151传递过来的值进行组合
assign value_variable_to_check_61[23:18] = value_variable_151_to_check_61;
assign enable_variable_to_check_61[3] = enable_variable_151_to_check_61;

// 拆分后校验节点61传递给变量节点202的值以及对变量节点202传递过来的值
wire [5:0] value_check_61_to_variable_202;
wire enable_check_61_to_variable_202;
wire [5:0] value_variable_202_to_check_61;
wire enable_variable_202_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_202 = value_check_61_to_variable[29:24];
assign enable_check_61_to_variable_202 = enable_check_61_to_variable[4];
// 对变量节点202传递过来的值进行组合
assign value_variable_to_check_61[29:24] = value_variable_202_to_check_61;
assign enable_variable_to_check_61[4] = enable_variable_202_to_check_61;

// 拆分后校验节点61传递给变量节点242的值以及对变量节点242传递过来的值
wire [5:0] value_check_61_to_variable_242;
wire enable_check_61_to_variable_242;
wire [5:0] value_variable_242_to_check_61;
wire enable_variable_242_to_check_61;
// 对校验节点61的输出值进行拆分
assign value_check_61_to_variable_242 = value_check_61_to_variable[35:30];
assign enable_check_61_to_variable_242 = enable_check_61_to_variable[5];
// 对变量节点242传递过来的值进行组合
assign value_variable_to_check_61[35:30] = value_variable_242_to_check_61;
assign enable_variable_to_check_61[5] = enable_variable_242_to_check_61;


// 校验节点62的接口
wire [35:0] value_variable_to_check_62;
wire [35:0] value_check_62_to_variable;
wire [5:0] enable_variable_to_check_62;
wire [5:0] enable_check_62_to_variable;

// 拆分后校验节点62传递给变量节点23的值以及对变量节点23传递过来的值
wire [5:0] value_check_62_to_variable_23;
wire enable_check_62_to_variable_23;
wire [5:0] value_variable_23_to_check_62;
wire enable_variable_23_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_23 = value_check_62_to_variable[5:0];
assign enable_check_62_to_variable_23 = enable_check_62_to_variable[0];
// 对变量节点23传递过来的值进行组合
assign value_variable_to_check_62[5:0] = value_variable_23_to_check_62;
assign enable_variable_to_check_62[0] = enable_variable_23_to_check_62;

// 拆分后校验节点62传递给变量节点57的值以及对变量节点57传递过来的值
wire [5:0] value_check_62_to_variable_57;
wire enable_check_62_to_variable_57;
wire [5:0] value_variable_57_to_check_62;
wire enable_variable_57_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_57 = value_check_62_to_variable[11:6];
assign enable_check_62_to_variable_57 = enable_check_62_to_variable[1];
// 对变量节点57传递过来的值进行组合
assign value_variable_to_check_62[11:6] = value_variable_57_to_check_62;
assign enable_variable_to_check_62[1] = enable_variable_57_to_check_62;

// 拆分后校验节点62传递给变量节点94的值以及对变量节点94传递过来的值
wire [5:0] value_check_62_to_variable_94;
wire enable_check_62_to_variable_94;
wire [5:0] value_variable_94_to_check_62;
wire enable_variable_94_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_94 = value_check_62_to_variable[17:12];
assign enable_check_62_to_variable_94 = enable_check_62_to_variable[2];
// 对变量节点94传递过来的值进行组合
assign value_variable_to_check_62[17:12] = value_variable_94_to_check_62;
assign enable_variable_to_check_62[2] = enable_variable_94_to_check_62;

// 拆分后校验节点62传递给变量节点132的值以及对变量节点132传递过来的值
wire [5:0] value_check_62_to_variable_132;
wire enable_check_62_to_variable_132;
wire [5:0] value_variable_132_to_check_62;
wire enable_variable_132_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_132 = value_check_62_to_variable[23:18];
assign enable_check_62_to_variable_132 = enable_check_62_to_variable[3];
// 对变量节点132传递过来的值进行组合
assign value_variable_to_check_62[23:18] = value_variable_132_to_check_62;
assign enable_variable_to_check_62[3] = enable_variable_132_to_check_62;

// 拆分后校验节点62传递给变量节点175的值以及对变量节点175传递过来的值
wire [5:0] value_check_62_to_variable_175;
wire enable_check_62_to_variable_175;
wire [5:0] value_variable_175_to_check_62;
wire enable_variable_175_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_175 = value_check_62_to_variable[29:24];
assign enable_check_62_to_variable_175 = enable_check_62_to_variable[4];
// 对变量节点175传递过来的值进行组合
assign value_variable_to_check_62[29:24] = value_variable_175_to_check_62;
assign enable_variable_to_check_62[4] = enable_variable_175_to_check_62;

// 拆分后校验节点62传递给变量节点248的值以及对变量节点248传递过来的值
wire [5:0] value_check_62_to_variable_248;
wire enable_check_62_to_variable_248;
wire [5:0] value_variable_248_to_check_62;
wire enable_variable_248_to_check_62;
// 对校验节点62的输出值进行拆分
assign value_check_62_to_variable_248 = value_check_62_to_variable[35:30];
assign enable_check_62_to_variable_248 = enable_check_62_to_variable[5];
// 对变量节点248传递过来的值进行组合
assign value_variable_to_check_62[35:30] = value_variable_248_to_check_62;
assign enable_variable_to_check_62[5] = enable_variable_248_to_check_62;


// 校验节点63的接口
wire [35:0] value_variable_to_check_63;
wire [35:0] value_check_63_to_variable;
wire [5:0] enable_variable_to_check_63;
wire [5:0] enable_check_63_to_variable;

// 拆分后校验节点63传递给变量节点22的值以及对变量节点22传递过来的值
wire [5:0] value_check_63_to_variable_22;
wire enable_check_63_to_variable_22;
wire [5:0] value_variable_22_to_check_63;
wire enable_variable_22_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_22 = value_check_63_to_variable[5:0];
assign enable_check_63_to_variable_22 = enable_check_63_to_variable[0];
// 对变量节点22传递过来的值进行组合
assign value_variable_to_check_63[5:0] = value_variable_22_to_check_63;
assign enable_variable_to_check_63[0] = enable_variable_22_to_check_63;

// 拆分后校验节点63传递给变量节点78的值以及对变量节点78传递过来的值
wire [5:0] value_check_63_to_variable_78;
wire enable_check_63_to_variable_78;
wire [5:0] value_variable_78_to_check_63;
wire enable_variable_78_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_78 = value_check_63_to_variable[11:6];
assign enable_check_63_to_variable_78 = enable_check_63_to_variable[1];
// 对变量节点78传递过来的值进行组合
assign value_variable_to_check_63[11:6] = value_variable_78_to_check_63;
assign enable_variable_to_check_63[1] = enable_variable_78_to_check_63;

// 拆分后校验节点63传递给变量节点113的值以及对变量节点113传递过来的值
wire [5:0] value_check_63_to_variable_113;
wire enable_check_63_to_variable_113;
wire [5:0] value_variable_113_to_check_63;
wire enable_variable_113_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_113 = value_check_63_to_variable[17:12];
assign enable_check_63_to_variable_113 = enable_check_63_to_variable[2];
// 对变量节点113传递过来的值进行组合
assign value_variable_to_check_63[17:12] = value_variable_113_to_check_63;
assign enable_variable_to_check_63[2] = enable_variable_113_to_check_63;

// 拆分后校验节点63传递给变量节点156的值以及对变量节点156传递过来的值
wire [5:0] value_check_63_to_variable_156;
wire enable_check_63_to_variable_156;
wire [5:0] value_variable_156_to_check_63;
wire enable_variable_156_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_156 = value_check_63_to_variable[23:18];
assign enable_check_63_to_variable_156 = enable_check_63_to_variable[3];
// 对变量节点156传递过来的值进行组合
assign value_variable_to_check_63[23:18] = value_variable_156_to_check_63;
assign enable_variable_to_check_63[3] = enable_variable_156_to_check_63;

// 拆分后校验节点63传递给变量节点207的值以及对变量节点207传递过来的值
wire [5:0] value_check_63_to_variable_207;
wire enable_check_63_to_variable_207;
wire [5:0] value_variable_207_to_check_63;
wire enable_variable_207_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_207 = value_check_63_to_variable[29:24];
assign enable_check_63_to_variable_207 = enable_check_63_to_variable[4];
// 对变量节点207传递过来的值进行组合
assign value_variable_to_check_63[29:24] = value_variable_207_to_check_63;
assign enable_variable_to_check_63[4] = enable_variable_207_to_check_63;

// 拆分后校验节点63传递给变量节点217的值以及对变量节点217传递过来的值
wire [5:0] value_check_63_to_variable_217;
wire enable_check_63_to_variable_217;
wire [5:0] value_variable_217_to_check_63;
wire enable_variable_217_to_check_63;
// 对校验节点63的输出值进行拆分
assign value_check_63_to_variable_217 = value_check_63_to_variable[35:30];
assign enable_check_63_to_variable_217 = enable_check_63_to_variable[5];
// 对变量节点217传递过来的值进行组合
assign value_variable_to_check_63[35:30] = value_variable_217_to_check_63;
assign enable_variable_to_check_63[5] = enable_variable_217_to_check_63;


// 校验节点64的接口
wire [35:0] value_variable_to_check_64;
wire [35:0] value_check_64_to_variable;
wire [5:0] enable_variable_to_check_64;
wire [5:0] enable_check_64_to_variable;

// 拆分后校验节点64传递给变量节点37的值以及对变量节点37传递过来的值
wire [5:0] value_check_64_to_variable_37;
wire enable_check_64_to_variable_37;
wire [5:0] value_variable_37_to_check_64;
wire enable_variable_37_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_37 = value_check_64_to_variable[5:0];
assign enable_check_64_to_variable_37 = enable_check_64_to_variable[0];
// 对变量节点37传递过来的值进行组合
assign value_variable_to_check_64[5:0] = value_variable_37_to_check_64;
assign enable_variable_to_check_64[0] = enable_variable_37_to_check_64;

// 拆分后校验节点64传递给变量节点79的值以及对变量节点79传递过来的值
wire [5:0] value_check_64_to_variable_79;
wire enable_check_64_to_variable_79;
wire [5:0] value_variable_79_to_check_64;
wire enable_variable_79_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_79 = value_check_64_to_variable[11:6];
assign enable_check_64_to_variable_79 = enable_check_64_to_variable[1];
// 对变量节点79传递过来的值进行组合
assign value_variable_to_check_64[11:6] = value_variable_79_to_check_64;
assign enable_variable_to_check_64[1] = enable_variable_79_to_check_64;

// 拆分后校验节点64传递给变量节点111的值以及对变量节点111传递过来的值
wire [5:0] value_check_64_to_variable_111;
wire enable_check_64_to_variable_111;
wire [5:0] value_variable_111_to_check_64;
wire enable_variable_111_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_111 = value_check_64_to_variable[17:12];
assign enable_check_64_to_variable_111 = enable_check_64_to_variable[2];
// 对变量节点111传递过来的值进行组合
assign value_variable_to_check_64[17:12] = value_variable_111_to_check_64;
assign enable_variable_to_check_64[2] = enable_variable_111_to_check_64;

// 拆分后校验节点64传递给变量节点127的值以及对变量节点127传递过来的值
wire [5:0] value_check_64_to_variable_127;
wire enable_check_64_to_variable_127;
wire [5:0] value_variable_127_to_check_64;
wire enable_variable_127_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_127 = value_check_64_to_variable[23:18];
assign enable_check_64_to_variable_127 = enable_check_64_to_variable[3];
// 对变量节点127传递过来的值进行组合
assign value_variable_to_check_64[23:18] = value_variable_127_to_check_64;
assign enable_variable_to_check_64[3] = enable_variable_127_to_check_64;

// 拆分后校验节点64传递给变量节点164的值以及对变量节点164传递过来的值
wire [5:0] value_check_64_to_variable_164;
wire enable_check_64_to_variable_164;
wire [5:0] value_variable_164_to_check_64;
wire enable_variable_164_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_164 = value_check_64_to_variable[29:24];
assign enable_check_64_to_variable_164 = enable_check_64_to_variable[4];
// 对变量节点164传递过来的值进行组合
assign value_variable_to_check_64[29:24] = value_variable_164_to_check_64;
assign enable_variable_to_check_64[4] = enable_variable_164_to_check_64;

// 拆分后校验节点64传递给变量节点239的值以及对变量节点239传递过来的值
wire [5:0] value_check_64_to_variable_239;
wire enable_check_64_to_variable_239;
wire [5:0] value_variable_239_to_check_64;
wire enable_variable_239_to_check_64;
// 对校验节点64的输出值进行拆分
assign value_check_64_to_variable_239 = value_check_64_to_variable[35:30];
assign enable_check_64_to_variable_239 = enable_check_64_to_variable[5];
// 对变量节点239传递过来的值进行组合
assign value_variable_to_check_64[35:30] = value_variable_239_to_check_64;
assign enable_variable_to_check_64[5] = enable_variable_239_to_check_64;


// 校验节点65的接口
wire [35:0] value_variable_to_check_65;
wire [35:0] value_check_65_to_variable;
wire [5:0] enable_variable_to_check_65;
wire [5:0] enable_check_65_to_variable;

// 拆分后校验节点65传递给变量节点24的值以及对变量节点24传递过来的值
wire [5:0] value_check_65_to_variable_24;
wire enable_check_65_to_variable_24;
wire [5:0] value_variable_24_to_check_65;
wire enable_variable_24_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_24 = value_check_65_to_variable[5:0];
assign enable_check_65_to_variable_24 = enable_check_65_to_variable[0];
// 对变量节点24传递过来的值进行组合
assign value_variable_to_check_65[5:0] = value_variable_24_to_check_65;
assign enable_variable_to_check_65[0] = enable_variable_24_to_check_65;

// 拆分后校验节点65传递给变量节点58的值以及对变量节点58传递过来的值
wire [5:0] value_check_65_to_variable_58;
wire enable_check_65_to_variable_58;
wire [5:0] value_variable_58_to_check_65;
wire enable_variable_58_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_58 = value_check_65_to_variable[11:6];
assign enable_check_65_to_variable_58 = enable_check_65_to_variable[1];
// 对变量节点58传递过来的值进行组合
assign value_variable_to_check_65[11:6] = value_variable_58_to_check_65;
assign enable_variable_to_check_65[1] = enable_variable_58_to_check_65;

// 拆分后校验节点65传递给变量节点114的值以及对变量节点114传递过来的值
wire [5:0] value_check_65_to_variable_114;
wire enable_check_65_to_variable_114;
wire [5:0] value_variable_114_to_check_65;
wire enable_variable_114_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_114 = value_check_65_to_variable[17:12];
assign enable_check_65_to_variable_114 = enable_check_65_to_variable[2];
// 对变量节点114传递过来的值进行组合
assign value_variable_to_check_65[17:12] = value_variable_114_to_check_65;
assign enable_variable_to_check_65[2] = enable_variable_114_to_check_65;

// 拆分后校验节点65传递给变量节点160的值以及对变量节点160传递过来的值
wire [5:0] value_check_65_to_variable_160;
wire enable_check_65_to_variable_160;
wire [5:0] value_variable_160_to_check_65;
wire enable_variable_160_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_160 = value_check_65_to_variable[23:18];
assign enable_check_65_to_variable_160 = enable_check_65_to_variable[3];
// 对变量节点160传递过来的值进行组合
assign value_variable_to_check_65[23:18] = value_variable_160_to_check_65;
assign enable_variable_to_check_65[3] = enable_variable_160_to_check_65;

// 拆分后校验节点65传递给变量节点197的值以及对变量节点197传递过来的值
wire [5:0] value_check_65_to_variable_197;
wire enable_check_65_to_variable_197;
wire [5:0] value_variable_197_to_check_65;
wire enable_variable_197_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_197 = value_check_65_to_variable[29:24];
assign enable_check_65_to_variable_197 = enable_check_65_to_variable[4];
// 对变量节点197传递过来的值进行组合
assign value_variable_to_check_65[29:24] = value_variable_197_to_check_65;
assign enable_variable_to_check_65[4] = enable_variable_197_to_check_65;

// 拆分后校验节点65传递给变量节点249的值以及对变量节点249传递过来的值
wire [5:0] value_check_65_to_variable_249;
wire enable_check_65_to_variable_249;
wire [5:0] value_variable_249_to_check_65;
wire enable_variable_249_to_check_65;
// 对校验节点65的输出值进行拆分
assign value_check_65_to_variable_249 = value_check_65_to_variable[35:30];
assign enable_check_65_to_variable_249 = enable_check_65_to_variable[5];
// 对变量节点249传递过来的值进行组合
assign value_variable_to_check_65[35:30] = value_variable_249_to_check_65;
assign enable_variable_to_check_65[5] = enable_variable_249_to_check_65;


// 校验节点66的接口
wire [35:0] value_variable_to_check_66;
wire [35:0] value_check_66_to_variable;
wire [5:0] enable_variable_to_check_66;
wire [5:0] enable_check_66_to_variable;

// 拆分后校验节点66传递给变量节点22的值以及对变量节点22传递过来的值
wire [5:0] value_check_66_to_variable_22;
wire enable_check_66_to_variable_22;
wire [5:0] value_variable_22_to_check_66;
wire enable_variable_22_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_22 = value_check_66_to_variable[5:0];
assign enable_check_66_to_variable_22 = enable_check_66_to_variable[0];
// 对变量节点22传递过来的值进行组合
assign value_variable_to_check_66[5:0] = value_variable_22_to_check_66;
assign enable_variable_to_check_66[0] = enable_variable_22_to_check_66;

// 拆分后校验节点66传递给变量节点80的值以及对变量节点80传递过来的值
wire [5:0] value_check_66_to_variable_80;
wire enable_check_66_to_variable_80;
wire [5:0] value_variable_80_to_check_66;
wire enable_variable_80_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_80 = value_check_66_to_variable[11:6];
assign enable_check_66_to_variable_80 = enable_check_66_to_variable[1];
// 对变量节点80传递过来的值进行组合
assign value_variable_to_check_66[11:6] = value_variable_80_to_check_66;
assign enable_variable_to_check_66[1] = enable_variable_80_to_check_66;

// 拆分后校验节点66传递给变量节点123的值以及对变量节点123传递过来的值
wire [5:0] value_check_66_to_variable_123;
wire enable_check_66_to_variable_123;
wire [5:0] value_variable_123_to_check_66;
wire enable_variable_123_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_123 = value_check_66_to_variable[17:12];
assign enable_check_66_to_variable_123 = enable_check_66_to_variable[2];
// 对变量节点123传递过来的值进行组合
assign value_variable_to_check_66[17:12] = value_variable_123_to_check_66;
assign enable_variable_to_check_66[2] = enable_variable_123_to_check_66;

// 拆分后校验节点66传递给变量节点130的值以及对变量节点130传递过来的值
wire [5:0] value_check_66_to_variable_130;
wire enable_check_66_to_variable_130;
wire [5:0] value_variable_130_to_check_66;
wire enable_variable_130_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_130 = value_check_66_to_variable[23:18];
assign enable_check_66_to_variable_130 = enable_check_66_to_variable[3];
// 对变量节点130传递过来的值进行组合
assign value_variable_to_check_66[23:18] = value_variable_130_to_check_66;
assign enable_variable_to_check_66[3] = enable_variable_130_to_check_66;

// 拆分后校验节点66传递给变量节点199的值以及对变量节点199传递过来的值
wire [5:0] value_check_66_to_variable_199;
wire enable_check_66_to_variable_199;
wire [5:0] value_variable_199_to_check_66;
wire enable_variable_199_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_199 = value_check_66_to_variable[29:24];
assign enable_check_66_to_variable_199 = enable_check_66_to_variable[4];
// 对变量节点199传递过来的值进行组合
assign value_variable_to_check_66[29:24] = value_variable_199_to_check_66;
assign enable_variable_to_check_66[4] = enable_variable_199_to_check_66;

// 拆分后校验节点66传递给变量节点248的值以及对变量节点248传递过来的值
wire [5:0] value_check_66_to_variable_248;
wire enable_check_66_to_variable_248;
wire [5:0] value_variable_248_to_check_66;
wire enable_variable_248_to_check_66;
// 对校验节点66的输出值进行拆分
assign value_check_66_to_variable_248 = value_check_66_to_variable[35:30];
assign enable_check_66_to_variable_248 = enable_check_66_to_variable[5];
// 对变量节点248传递过来的值进行组合
assign value_variable_to_check_66[35:30] = value_variable_248_to_check_66;
assign enable_variable_to_check_66[5] = enable_variable_248_to_check_66;


// 校验节点67的接口
wire [35:0] value_variable_to_check_67;
wire [35:0] value_check_67_to_variable;
wire [5:0] enable_variable_to_check_67;
wire [5:0] enable_check_67_to_variable;

// 拆分后校验节点67传递给变量节点31的值以及对变量节点31传递过来的值
wire [5:0] value_check_67_to_variable_31;
wire enable_check_67_to_variable_31;
wire [5:0] value_variable_31_to_check_67;
wire enable_variable_31_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_31 = value_check_67_to_variable[5:0];
assign enable_check_67_to_variable_31 = enable_check_67_to_variable[0];
// 对变量节点31传递过来的值进行组合
assign value_variable_to_check_67[5:0] = value_variable_31_to_check_67;
assign enable_variable_to_check_67[0] = enable_variable_31_to_check_67;

// 拆分后校验节点67传递给变量节点81的值以及对变量节点81传递过来的值
wire [5:0] value_check_67_to_variable_81;
wire enable_check_67_to_variable_81;
wire [5:0] value_variable_81_to_check_67;
wire enable_variable_81_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_81 = value_check_67_to_variable[11:6];
assign enable_check_67_to_variable_81 = enable_check_67_to_variable[1];
// 对变量节点81传递过来的值进行组合
assign value_variable_to_check_67[11:6] = value_variable_81_to_check_67;
assign enable_variable_to_check_67[1] = enable_variable_81_to_check_67;

// 拆分后校验节点67传递给变量节点91的值以及对变量节点91传递过来的值
wire [5:0] value_check_67_to_variable_91;
wire enable_check_67_to_variable_91;
wire [5:0] value_variable_91_to_check_67;
wire enable_variable_91_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_91 = value_check_67_to_variable[17:12];
assign enable_check_67_to_variable_91 = enable_check_67_to_variable[2];
// 对变量节点91传递过来的值进行组合
assign value_variable_to_check_67[17:12] = value_variable_91_to_check_67;
assign enable_variable_to_check_67[2] = enable_variable_91_to_check_67;

// 拆分后校验节点67传递给变量节点164的值以及对变量节点164传递过来的值
wire [5:0] value_check_67_to_variable_164;
wire enable_check_67_to_variable_164;
wire [5:0] value_variable_164_to_check_67;
wire enable_variable_164_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_164 = value_check_67_to_variable[23:18];
assign enable_check_67_to_variable_164 = enable_check_67_to_variable[3];
// 对变量节点164传递过来的值进行组合
assign value_variable_to_check_67[23:18] = value_variable_164_to_check_67;
assign enable_variable_to_check_67[3] = enable_variable_164_to_check_67;

// 拆分后校验节点67传递给变量节点180的值以及对变量节点180传递过来的值
wire [5:0] value_check_67_to_variable_180;
wire enable_check_67_to_variable_180;
wire [5:0] value_variable_180_to_check_67;
wire enable_variable_180_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_180 = value_check_67_to_variable[29:24];
assign enable_check_67_to_variable_180 = enable_check_67_to_variable[4];
// 对变量节点180传递过来的值进行组合
assign value_variable_to_check_67[29:24] = value_variable_180_to_check_67;
assign enable_variable_to_check_67[4] = enable_variable_180_to_check_67;

// 拆分后校验节点67传递给变量节点223的值以及对变量节点223传递过来的值
wire [5:0] value_check_67_to_variable_223;
wire enable_check_67_to_variable_223;
wire [5:0] value_variable_223_to_check_67;
wire enable_variable_223_to_check_67;
// 对校验节点67的输出值进行拆分
assign value_check_67_to_variable_223 = value_check_67_to_variable[35:30];
assign enable_check_67_to_variable_223 = enable_check_67_to_variable[5];
// 对变量节点223传递过来的值进行组合
assign value_variable_to_check_67[35:30] = value_variable_223_to_check_67;
assign enable_variable_to_check_67[5] = enable_variable_223_to_check_67;


// 校验节点68的接口
wire [35:0] value_variable_to_check_68;
wire [35:0] value_check_68_to_variable;
wire [5:0] enable_variable_to_check_68;
wire [5:0] enable_check_68_to_variable;

// 拆分后校验节点68传递给变量节点38的值以及对变量节点38传递过来的值
wire [5:0] value_check_68_to_variable_38;
wire enable_check_68_to_variable_38;
wire [5:0] value_variable_38_to_check_68;
wire enable_variable_38_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_38 = value_check_68_to_variable[5:0];
assign enable_check_68_to_variable_38 = enable_check_68_to_variable[0];
// 对变量节点38传递过来的值进行组合
assign value_variable_to_check_68[5:0] = value_variable_38_to_check_68;
assign enable_variable_to_check_68[0] = enable_variable_38_to_check_68;

// 拆分后校验节点68传递给变量节点78的值以及对变量节点78传递过来的值
wire [5:0] value_check_68_to_variable_78;
wire enable_check_68_to_variable_78;
wire [5:0] value_variable_78_to_check_68;
wire enable_variable_78_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_78 = value_check_68_to_variable[11:6];
assign enable_check_68_to_variable_78 = enable_check_68_to_variable[1];
// 对变量节点78传递过来的值进行组合
assign value_variable_to_check_68[11:6] = value_variable_78_to_check_68;
assign enable_variable_to_check_68[1] = enable_variable_78_to_check_68;

// 拆分后校验节点68传递给变量节点88的值以及对变量节点88传递过来的值
wire [5:0] value_check_68_to_variable_88;
wire enable_check_68_to_variable_88;
wire [5:0] value_variable_88_to_check_68;
wire enable_variable_88_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_88 = value_check_68_to_variable[17:12];
assign enable_check_68_to_variable_88 = enable_check_68_to_variable[2];
// 对变量节点88传递过来的值进行组合
assign value_variable_to_check_68[17:12] = value_variable_88_to_check_68;
assign enable_variable_to_check_68[2] = enable_variable_88_to_check_68;

// 拆分后校验节点68传递给变量节点160的值以及对变量节点160传递过来的值
wire [5:0] value_check_68_to_variable_160;
wire enable_check_68_to_variable_160;
wire [5:0] value_variable_160_to_check_68;
wire enable_variable_160_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_160 = value_check_68_to_variable[23:18];
assign enable_check_68_to_variable_160 = enable_check_68_to_variable[3];
// 对变量节点160传递过来的值进行组合
assign value_variable_to_check_68[23:18] = value_variable_160_to_check_68;
assign enable_variable_to_check_68[3] = enable_variable_160_to_check_68;

// 拆分后校验节点68传递给变量节点208的值以及对变量节点208传递过来的值
wire [5:0] value_check_68_to_variable_208;
wire enable_check_68_to_variable_208;
wire [5:0] value_variable_208_to_check_68;
wire enable_variable_208_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_208 = value_check_68_to_variable[29:24];
assign enable_check_68_to_variable_208 = enable_check_68_to_variable[4];
// 对变量节点208传递过来的值进行组合
assign value_variable_to_check_68[29:24] = value_variable_208_to_check_68;
assign enable_variable_to_check_68[4] = enable_variable_208_to_check_68;

// 拆分后校验节点68传递给变量节点250的值以及对变量节点250传递过来的值
wire [5:0] value_check_68_to_variable_250;
wire enable_check_68_to_variable_250;
wire [5:0] value_variable_250_to_check_68;
wire enable_variable_250_to_check_68;
// 对校验节点68的输出值进行拆分
assign value_check_68_to_variable_250 = value_check_68_to_variable[35:30];
assign enable_check_68_to_variable_250 = enable_check_68_to_variable[5];
// 对变量节点250传递过来的值进行组合
assign value_variable_to_check_68[35:30] = value_variable_250_to_check_68;
assign enable_variable_to_check_68[5] = enable_variable_250_to_check_68;


// 校验节点69的接口
wire [35:0] value_variable_to_check_69;
wire [35:0] value_check_69_to_variable;
wire [5:0] enable_variable_to_check_69;
wire [5:0] enable_check_69_to_variable;

// 拆分后校验节点69传递给变量节点38的值以及对变量节点38传递过来的值
wire [5:0] value_check_69_to_variable_38;
wire enable_check_69_to_variable_38;
wire [5:0] value_variable_38_to_check_69;
wire enable_variable_38_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_38 = value_check_69_to_variable[5:0];
assign enable_check_69_to_variable_38 = enable_check_69_to_variable[0];
// 对变量节点38传递过来的值进行组合
assign value_variable_to_check_69[5:0] = value_variable_38_to_check_69;
assign enable_variable_to_check_69[0] = enable_variable_38_to_check_69;

// 拆分后校验节点69传递给变量节点48的值以及对变量节点48传递过来的值
wire [5:0] value_check_69_to_variable_48;
wire enable_check_69_to_variable_48;
wire [5:0] value_variable_48_to_check_69;
wire enable_variable_48_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_48 = value_check_69_to_variable[11:6];
assign enable_check_69_to_variable_48 = enable_check_69_to_variable[1];
// 对变量节点48传递过来的值进行组合
assign value_variable_to_check_69[11:6] = value_variable_48_to_check_69;
assign enable_variable_to_check_69[1] = enable_variable_48_to_check_69;

// 拆分后校验节点69传递给变量节点110的值以及对变量节点110传递过来的值
wire [5:0] value_check_69_to_variable_110;
wire enable_check_69_to_variable_110;
wire [5:0] value_variable_110_to_check_69;
wire enable_variable_110_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_110 = value_check_69_to_variable[17:12];
assign enable_check_69_to_variable_110 = enable_check_69_to_variable[2];
// 对变量节点110传递过来的值进行组合
assign value_variable_to_check_69[17:12] = value_variable_110_to_check_69;
assign enable_variable_to_check_69[2] = enable_variable_110_to_check_69;

// 拆分后校验节点69传递给变量节点139的值以及对变量节点139传递过来的值
wire [5:0] value_check_69_to_variable_139;
wire enable_check_69_to_variable_139;
wire [5:0] value_variable_139_to_check_69;
wire enable_variable_139_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_139 = value_check_69_to_variable[23:18];
assign enable_check_69_to_variable_139 = enable_check_69_to_variable[3];
// 对变量节点139传递过来的值进行组合
assign value_variable_to_check_69[23:18] = value_variable_139_to_check_69;
assign enable_variable_to_check_69[3] = enable_variable_139_to_check_69;

// 拆分后校验节点69传递给变量节点177的值以及对变量节点177传递过来的值
wire [5:0] value_check_69_to_variable_177;
wire enable_check_69_to_variable_177;
wire [5:0] value_variable_177_to_check_69;
wire enable_variable_177_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_177 = value_check_69_to_variable[29:24];
assign enable_check_69_to_variable_177 = enable_check_69_to_variable[4];
// 对变量节点177传递过来的值进行组合
assign value_variable_to_check_69[29:24] = value_variable_177_to_check_69;
assign enable_variable_to_check_69[4] = enable_variable_177_to_check_69;

// 拆分后校验节点69传递给变量节点212的值以及对变量节点212传递过来的值
wire [5:0] value_check_69_to_variable_212;
wire enable_check_69_to_variable_212;
wire [5:0] value_variable_212_to_check_69;
wire enable_variable_212_to_check_69;
// 对校验节点69的输出值进行拆分
assign value_check_69_to_variable_212 = value_check_69_to_variable[35:30];
assign enable_check_69_to_variable_212 = enable_check_69_to_variable[5];
// 对变量节点212传递过来的值进行组合
assign value_variable_to_check_69[35:30] = value_variable_212_to_check_69;
assign enable_variable_to_check_69[5] = enable_variable_212_to_check_69;


// 校验节点70的接口
wire [35:0] value_variable_to_check_70;
wire [35:0] value_check_70_to_variable;
wire [5:0] enable_variable_to_check_70;
wire [5:0] enable_check_70_to_variable;

// 拆分后校验节点70传递给变量节点39的值以及对变量节点39传递过来的值
wire [5:0] value_check_70_to_variable_39;
wire enable_check_70_to_variable_39;
wire [5:0] value_variable_39_to_check_70;
wire enable_variable_39_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_39 = value_check_70_to_variable[5:0];
assign enable_check_70_to_variable_39 = enable_check_70_to_variable[0];
// 对变量节点39传递过来的值进行组合
assign value_variable_to_check_70[5:0] = value_variable_39_to_check_70;
assign enable_variable_to_check_70[0] = enable_variable_39_to_check_70;

// 拆分后校验节点70传递给变量节点53的值以及对变量节点53传递过来的值
wire [5:0] value_check_70_to_variable_53;
wire enable_check_70_to_variable_53;
wire [5:0] value_variable_53_to_check_70;
wire enable_variable_53_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_53 = value_check_70_to_variable[11:6];
assign enable_check_70_to_variable_53 = enable_check_70_to_variable[1];
// 对变量节点53传递过来的值进行组合
assign value_variable_to_check_70[11:6] = value_variable_53_to_check_70;
assign enable_variable_to_check_70[1] = enable_variable_53_to_check_70;

// 拆分后校验节点70传递给变量节点124的值以及对变量节点124传递过来的值
wire [5:0] value_check_70_to_variable_124;
wire enable_check_70_to_variable_124;
wire [5:0] value_variable_124_to_check_70;
wire enable_variable_124_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_124 = value_check_70_to_variable[17:12];
assign enable_check_70_to_variable_124 = enable_check_70_to_variable[2];
// 对变量节点124传递过来的值进行组合
assign value_variable_to_check_70[17:12] = value_variable_124_to_check_70;
assign enable_variable_to_check_70[2] = enable_variable_124_to_check_70;

// 拆分后校验节点70传递给变量节点150的值以及对变量节点150传递过来的值
wire [5:0] value_check_70_to_variable_150;
wire enable_check_70_to_variable_150;
wire [5:0] value_variable_150_to_check_70;
wire enable_variable_150_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_150 = value_check_70_to_variable[23:18];
assign enable_check_70_to_variable_150 = enable_check_70_to_variable[3];
// 对变量节点150传递过来的值进行组合
assign value_variable_to_check_70[23:18] = value_variable_150_to_check_70;
assign enable_variable_to_check_70[3] = enable_variable_150_to_check_70;

// 拆分后校验节点70传递给变量节点197的值以及对变量节点197传递过来的值
wire [5:0] value_check_70_to_variable_197;
wire enable_check_70_to_variable_197;
wire [5:0] value_variable_197_to_check_70;
wire enable_variable_197_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_197 = value_check_70_to_variable[29:24];
assign enable_check_70_to_variable_197 = enable_check_70_to_variable[4];
// 对变量节点197传递过来的值进行组合
assign value_variable_to_check_70[29:24] = value_variable_197_to_check_70;
assign enable_variable_to_check_70[4] = enable_variable_197_to_check_70;

// 拆分后校验节点70传递给变量节点251的值以及对变量节点251传递过来的值
wire [5:0] value_check_70_to_variable_251;
wire enable_check_70_to_variable_251;
wire [5:0] value_variable_251_to_check_70;
wire enable_variable_251_to_check_70;
// 对校验节点70的输出值进行拆分
assign value_check_70_to_variable_251 = value_check_70_to_variable[35:30];
assign enable_check_70_to_variable_251 = enable_check_70_to_variable[5];
// 对变量节点251传递过来的值进行组合
assign value_variable_to_check_70[35:30] = value_variable_251_to_check_70;
assign enable_variable_to_check_70[5] = enable_variable_251_to_check_70;


// 校验节点71的接口
wire [35:0] value_variable_to_check_71;
wire [35:0] value_check_71_to_variable;
wire [5:0] enable_variable_to_check_71;
wire [5:0] enable_check_71_to_variable;

// 拆分后校验节点71传递给变量节点40的值以及对变量节点40传递过来的值
wire [5:0] value_check_71_to_variable_40;
wire enable_check_71_to_variable_40;
wire [5:0] value_variable_40_to_check_71;
wire enable_variable_40_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_40 = value_check_71_to_variable[5:0];
assign enable_check_71_to_variable_40 = enable_check_71_to_variable[0];
// 对变量节点40传递过来的值进行组合
assign value_variable_to_check_71[5:0] = value_variable_40_to_check_71;
assign enable_variable_to_check_71[0] = enable_variable_40_to_check_71;

// 拆分后校验节点71传递给变量节点61的值以及对变量节点61传递过来的值
wire [5:0] value_check_71_to_variable_61;
wire enable_check_71_to_variable_61;
wire [5:0] value_variable_61_to_check_71;
wire enable_variable_61_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_61 = value_check_71_to_variable[11:6];
assign enable_check_71_to_variable_61 = enable_check_71_to_variable[1];
// 对变量节点61传递过来的值进行组合
assign value_variable_to_check_71[11:6] = value_variable_61_to_check_71;
assign enable_variable_to_check_71[1] = enable_variable_61_to_check_71;

// 拆分后校验节点71传递给变量节点110的值以及对变量节点110传递过来的值
wire [5:0] value_check_71_to_variable_110;
wire enable_check_71_to_variable_110;
wire [5:0] value_variable_110_to_check_71;
wire enable_variable_110_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_110 = value_check_71_to_variable[17:12];
assign enable_check_71_to_variable_110 = enable_check_71_to_variable[2];
// 对变量节点110传递过来的值进行组合
assign value_variable_to_check_71[17:12] = value_variable_110_to_check_71;
assign enable_variable_to_check_71[2] = enable_variable_110_to_check_71;

// 拆分后校验节点71传递给变量节点158的值以及对变量节点158传递过来的值
wire [5:0] value_check_71_to_variable_158;
wire enable_check_71_to_variable_158;
wire [5:0] value_variable_158_to_check_71;
wire enable_variable_158_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_158 = value_check_71_to_variable[23:18];
assign enable_check_71_to_variable_158 = enable_check_71_to_variable[3];
// 对变量节点158传递过来的值进行组合
assign value_variable_to_check_71[23:18] = value_variable_158_to_check_71;
assign enable_variable_to_check_71[3] = enable_variable_158_to_check_71;

// 拆分后校验节点71传递给变量节点191的值以及对变量节点191传递过来的值
wire [5:0] value_check_71_to_variable_191;
wire enable_check_71_to_variable_191;
wire [5:0] value_variable_191_to_check_71;
wire enable_variable_191_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_191 = value_check_71_to_variable[29:24];
assign enable_check_71_to_variable_191 = enable_check_71_to_variable[4];
// 对变量节点191传递过来的值进行组合
assign value_variable_to_check_71[29:24] = value_variable_191_to_check_71;
assign enable_variable_to_check_71[4] = enable_variable_191_to_check_71;

// 拆分后校验节点71传递给变量节点227的值以及对变量节点227传递过来的值
wire [5:0] value_check_71_to_variable_227;
wire enable_check_71_to_variable_227;
wire [5:0] value_variable_227_to_check_71;
wire enable_variable_227_to_check_71;
// 对校验节点71的输出值进行拆分
assign value_check_71_to_variable_227 = value_check_71_to_variable[35:30];
assign enable_check_71_to_variable_227 = enable_check_71_to_variable[5];
// 对变量节点227传递过来的值进行组合
assign value_variable_to_check_71[35:30] = value_variable_227_to_check_71;
assign enable_variable_to_check_71[5] = enable_variable_227_to_check_71;


// 校验节点72的接口
wire [35:0] value_variable_to_check_72;
wire [35:0] value_check_72_to_variable;
wire [5:0] enable_variable_to_check_72;
wire [5:0] enable_check_72_to_variable;

// 拆分后校验节点72传递给变量节点15的值以及对变量节点15传递过来的值
wire [5:0] value_check_72_to_variable_15;
wire enable_check_72_to_variable_15;
wire [5:0] value_variable_15_to_check_72;
wire enable_variable_15_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_15 = value_check_72_to_variable[5:0];
assign enable_check_72_to_variable_15 = enable_check_72_to_variable[0];
// 对变量节点15传递过来的值进行组合
assign value_variable_to_check_72[5:0] = value_variable_15_to_check_72;
assign enable_variable_to_check_72[0] = enable_variable_15_to_check_72;

// 拆分后校验节点72传递给变量节点44的值以及对变量节点44传递过来的值
wire [5:0] value_check_72_to_variable_44;
wire enable_check_72_to_variable_44;
wire [5:0] value_variable_44_to_check_72;
wire enable_variable_44_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_44 = value_check_72_to_variable[11:6];
assign enable_check_72_to_variable_44 = enable_check_72_to_variable[1];
// 对变量节点44传递过来的值进行组合
assign value_variable_to_check_72[11:6] = value_variable_44_to_check_72;
assign enable_variable_to_check_72[1] = enable_variable_44_to_check_72;

// 拆分后校验节点72传递给变量节点86的值以及对变量节点86传递过来的值
wire [5:0] value_check_72_to_variable_86;
wire enable_check_72_to_variable_86;
wire [5:0] value_variable_86_to_check_72;
wire enable_variable_86_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_86 = value_check_72_to_variable[17:12];
assign enable_check_72_to_variable_86 = enable_check_72_to_variable[2];
// 对变量节点86传递过来的值进行组合
assign value_variable_to_check_72[17:12] = value_variable_86_to_check_72;
assign enable_variable_to_check_72[2] = enable_variable_86_to_check_72;

// 拆分后校验节点72传递给变量节点165的值以及对变量节点165传递过来的值
wire [5:0] value_check_72_to_variable_165;
wire enable_check_72_to_variable_165;
wire [5:0] value_variable_165_to_check_72;
wire enable_variable_165_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_165 = value_check_72_to_variable[23:18];
assign enable_check_72_to_variable_165 = enable_check_72_to_variable[3];
// 对变量节点165传递过来的值进行组合
assign value_variable_to_check_72[23:18] = value_variable_165_to_check_72;
assign enable_variable_to_check_72[3] = enable_variable_165_to_check_72;

// 拆分后校验节点72传递给变量节点206的值以及对变量节点206传递过来的值
wire [5:0] value_check_72_to_variable_206;
wire enable_check_72_to_variable_206;
wire [5:0] value_variable_206_to_check_72;
wire enable_variable_206_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_206 = value_check_72_to_variable[29:24];
assign enable_check_72_to_variable_206 = enable_check_72_to_variable[4];
// 对变量节点206传递过来的值进行组合
assign value_variable_to_check_72[29:24] = value_variable_206_to_check_72;
assign enable_variable_to_check_72[4] = enable_variable_206_to_check_72;

// 拆分后校验节点72传递给变量节点252的值以及对变量节点252传递过来的值
wire [5:0] value_check_72_to_variable_252;
wire enable_check_72_to_variable_252;
wire [5:0] value_variable_252_to_check_72;
wire enable_variable_252_to_check_72;
// 对校验节点72的输出值进行拆分
assign value_check_72_to_variable_252 = value_check_72_to_variable[35:30];
assign enable_check_72_to_variable_252 = enable_check_72_to_variable[5];
// 对变量节点252传递过来的值进行组合
assign value_variable_to_check_72[35:30] = value_variable_252_to_check_72;
assign enable_variable_to_check_72[5] = enable_variable_252_to_check_72;


// 校验节点73的接口
wire [35:0] value_variable_to_check_73;
wire [35:0] value_check_73_to_variable;
wire [5:0] enable_variable_to_check_73;
wire [5:0] enable_check_73_to_variable;

// 拆分后校验节点73传递给变量节点6的值以及对变量节点6传递过来的值
wire [5:0] value_check_73_to_variable_6;
wire enable_check_73_to_variable_6;
wire [5:0] value_variable_6_to_check_73;
wire enable_variable_6_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_6 = value_check_73_to_variable[5:0];
assign enable_check_73_to_variable_6 = enable_check_73_to_variable[0];
// 对变量节点6传递过来的值进行组合
assign value_variable_to_check_73[5:0] = value_variable_6_to_check_73;
assign enable_variable_to_check_73[0] = enable_variable_6_to_check_73;

// 拆分后校验节点73传递给变量节点77的值以及对变量节点77传递过来的值
wire [5:0] value_check_73_to_variable_77;
wire enable_check_73_to_variable_77;
wire [5:0] value_variable_77_to_check_73;
wire enable_variable_77_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_77 = value_check_73_to_variable[11:6];
assign enable_check_73_to_variable_77 = enable_check_73_to_variable[1];
// 对变量节点77传递过来的值进行组合
assign value_variable_to_check_73[11:6] = value_variable_77_to_check_73;
assign enable_variable_to_check_73[1] = enable_variable_77_to_check_73;

// 拆分后校验节点73传递给变量节点96的值以及对变量节点96传递过来的值
wire [5:0] value_check_73_to_variable_96;
wire enable_check_73_to_variable_96;
wire [5:0] value_variable_96_to_check_73;
wire enable_variable_96_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_96 = value_check_73_to_variable[17:12];
assign enable_check_73_to_variable_96 = enable_check_73_to_variable[2];
// 对变量节点96传递过来的值进行组合
assign value_variable_to_check_73[17:12] = value_variable_96_to_check_73;
assign enable_variable_to_check_73[2] = enable_variable_96_to_check_73;

// 拆分后校验节点73传递给变量节点156的值以及对变量节点156传递过来的值
wire [5:0] value_check_73_to_variable_156;
wire enable_check_73_to_variable_156;
wire [5:0] value_variable_156_to_check_73;
wire enable_variable_156_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_156 = value_check_73_to_variable[23:18];
assign enable_check_73_to_variable_156 = enable_check_73_to_variable[3];
// 对变量节点156传递过来的值进行组合
assign value_variable_to_check_73[23:18] = value_variable_156_to_check_73;
assign enable_variable_to_check_73[3] = enable_variable_156_to_check_73;

// 拆分后校验节点73传递给变量节点209的值以及对变量节点209传递过来的值
wire [5:0] value_check_73_to_variable_209;
wire enable_check_73_to_variable_209;
wire [5:0] value_variable_209_to_check_73;
wire enable_variable_209_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_209 = value_check_73_to_variable[29:24];
assign enable_check_73_to_variable_209 = enable_check_73_to_variable[4];
// 对变量节点209传递过来的值进行组合
assign value_variable_to_check_73[29:24] = value_variable_209_to_check_73;
assign enable_variable_to_check_73[4] = enable_variable_209_to_check_73;

// 拆分后校验节点73传递给变量节点216的值以及对变量节点216传递过来的值
wire [5:0] value_check_73_to_variable_216;
wire enable_check_73_to_variable_216;
wire [5:0] value_variable_216_to_check_73;
wire enable_variable_216_to_check_73;
// 对校验节点73的输出值进行拆分
assign value_check_73_to_variable_216 = value_check_73_to_variable[35:30];
assign enable_check_73_to_variable_216 = enable_check_73_to_variable[5];
// 对变量节点216传递过来的值进行组合
assign value_variable_to_check_73[35:30] = value_variable_216_to_check_73;
assign enable_variable_to_check_73[5] = enable_variable_216_to_check_73;


// 校验节点74的接口
wire [35:0] value_variable_to_check_74;
wire [35:0] value_check_74_to_variable;
wire [5:0] enable_variable_to_check_74;
wire [5:0] enable_check_74_to_variable;

// 拆分后校验节点74传递给变量节点3的值以及对变量节点3传递过来的值
wire [5:0] value_check_74_to_variable_3;
wire enable_check_74_to_variable_3;
wire [5:0] value_variable_3_to_check_74;
wire enable_variable_3_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_3 = value_check_74_to_variable[5:0];
assign enable_check_74_to_variable_3 = enable_check_74_to_variable[0];
// 对变量节点3传递过来的值进行组合
assign value_variable_to_check_74[5:0] = value_variable_3_to_check_74;
assign enable_variable_to_check_74[0] = enable_variable_3_to_check_74;

// 拆分后校验节点74传递给变量节点48的值以及对变量节点48传递过来的值
wire [5:0] value_check_74_to_variable_48;
wire enable_check_74_to_variable_48;
wire [5:0] value_variable_48_to_check_74;
wire enable_variable_48_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_48 = value_check_74_to_variable[11:6];
assign enable_check_74_to_variable_48 = enable_check_74_to_variable[1];
// 对变量节点48传递过来的值进行组合
assign value_variable_to_check_74[11:6] = value_variable_48_to_check_74;
assign enable_variable_to_check_74[1] = enable_variable_48_to_check_74;

// 拆分后校验节点74传递给变量节点125的值以及对变量节点125传递过来的值
wire [5:0] value_check_74_to_variable_125;
wire enable_check_74_to_variable_125;
wire [5:0] value_variable_125_to_check_74;
wire enable_variable_125_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_125 = value_check_74_to_variable[17:12];
assign enable_check_74_to_variable_125 = enable_check_74_to_variable[2];
// 对变量节点125传递过来的值进行组合
assign value_variable_to_check_74[17:12] = value_variable_125_to_check_74;
assign enable_variable_to_check_74[2] = enable_variable_125_to_check_74;

// 拆分后校验节点74传递给变量节点130的值以及对变量节点130传递过来的值
wire [5:0] value_check_74_to_variable_130;
wire enable_check_74_to_variable_130;
wire [5:0] value_variable_130_to_check_74;
wire enable_variable_130_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_130 = value_check_74_to_variable[23:18];
assign enable_check_74_to_variable_130 = enable_check_74_to_variable[3];
// 对变量节点130传递过来的值进行组合
assign value_variable_to_check_74[23:18] = value_variable_130_to_check_74;
assign enable_variable_to_check_74[3] = enable_variable_130_to_check_74;

// 拆分后校验节点74传递给变量节点188的值以及对变量节点188传递过来的值
wire [5:0] value_check_74_to_variable_188;
wire enable_check_74_to_variable_188;
wire [5:0] value_variable_188_to_check_74;
wire enable_variable_188_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_188 = value_check_74_to_variable[29:24];
assign enable_check_74_to_variable_188 = enable_check_74_to_variable[4];
// 对变量节点188传递过来的值进行组合
assign value_variable_to_check_74[29:24] = value_variable_188_to_check_74;
assign enable_variable_to_check_74[4] = enable_variable_188_to_check_74;

// 拆分后校验节点74传递给变量节点249的值以及对变量节点249传递过来的值
wire [5:0] value_check_74_to_variable_249;
wire enable_check_74_to_variable_249;
wire [5:0] value_variable_249_to_check_74;
wire enable_variable_249_to_check_74;
// 对校验节点74的输出值进行拆分
assign value_check_74_to_variable_249 = value_check_74_to_variable[35:30];
assign enable_check_74_to_variable_249 = enable_check_74_to_variable[5];
// 对变量节点249传递过来的值进行组合
assign value_variable_to_check_74[35:30] = value_variable_249_to_check_74;
assign enable_variable_to_check_74[5] = enable_variable_249_to_check_74;


// 校验节点75的接口
wire [35:0] value_variable_to_check_75;
wire [35:0] value_check_75_to_variable;
wire [5:0] enable_variable_to_check_75;
wire [5:0] enable_check_75_to_variable;

// 拆分后校验节点75传递给变量节点26的值以及对变量节点26传递过来的值
wire [5:0] value_check_75_to_variable_26;
wire enable_check_75_to_variable_26;
wire [5:0] value_variable_26_to_check_75;
wire enable_variable_26_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_26 = value_check_75_to_variable[5:0];
assign enable_check_75_to_variable_26 = enable_check_75_to_variable[0];
// 对变量节点26传递过来的值进行组合
assign value_variable_to_check_75[5:0] = value_variable_26_to_check_75;
assign enable_variable_to_check_75[0] = enable_variable_26_to_check_75;

// 拆分后校验节点75传递给变量节点81的值以及对变量节点81传递过来的值
wire [5:0] value_check_75_to_variable_81;
wire enable_check_75_to_variable_81;
wire [5:0] value_variable_81_to_check_75;
wire enable_variable_81_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_81 = value_check_75_to_variable[11:6];
assign enable_check_75_to_variable_81 = enable_check_75_to_variable[1];
// 对变量节点81传递过来的值进行组合
assign value_variable_to_check_75[11:6] = value_variable_81_to_check_75;
assign enable_variable_to_check_75[1] = enable_variable_81_to_check_75;

// 拆分后校验节点75传递给变量节点103的值以及对变量节点103传递过来的值
wire [5:0] value_check_75_to_variable_103;
wire enable_check_75_to_variable_103;
wire [5:0] value_variable_103_to_check_75;
wire enable_variable_103_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_103 = value_check_75_to_variable[17:12];
assign enable_check_75_to_variable_103 = enable_check_75_to_variable[2];
// 对变量节点103传递过来的值进行组合
assign value_variable_to_check_75[17:12] = value_variable_103_to_check_75;
assign enable_variable_to_check_75[2] = enable_variable_103_to_check_75;

// 拆分后校验节点75传递给变量节点141的值以及对变量节点141传递过来的值
wire [5:0] value_check_75_to_variable_141;
wire enable_check_75_to_variable_141;
wire [5:0] value_variable_141_to_check_75;
wire enable_variable_141_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_141 = value_check_75_to_variable[23:18];
assign enable_check_75_to_variable_141 = enable_check_75_to_variable[3];
// 对变量节点141传递过来的值进行组合
assign value_variable_to_check_75[23:18] = value_variable_141_to_check_75;
assign enable_variable_to_check_75[3] = enable_variable_141_to_check_75;

// 拆分后校验节点75传递给变量节点200的值以及对变量节点200传递过来的值
wire [5:0] value_check_75_to_variable_200;
wire enable_check_75_to_variable_200;
wire [5:0] value_variable_200_to_check_75;
wire enable_variable_200_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_200 = value_check_75_to_variable[29:24];
assign enable_check_75_to_variable_200 = enable_check_75_to_variable[4];
// 对变量节点200传递过来的值进行组合
assign value_variable_to_check_75[29:24] = value_variable_200_to_check_75;
assign enable_variable_to_check_75[4] = enable_variable_200_to_check_75;

// 拆分后校验节点75传递给变量节点234的值以及对变量节点234传递过来的值
wire [5:0] value_check_75_to_variable_234;
wire enable_check_75_to_variable_234;
wire [5:0] value_variable_234_to_check_75;
wire enable_variable_234_to_check_75;
// 对校验节点75的输出值进行拆分
assign value_check_75_to_variable_234 = value_check_75_to_variable[35:30];
assign enable_check_75_to_variable_234 = enable_check_75_to_variable[5];
// 对变量节点234传递过来的值进行组合
assign value_variable_to_check_75[35:30] = value_variable_234_to_check_75;
assign enable_variable_to_check_75[5] = enable_variable_234_to_check_75;


// 校验节点76的接口
wire [35:0] value_variable_to_check_76;
wire [35:0] value_check_76_to_variable;
wire [5:0] enable_variable_to_check_76;
wire [5:0] enable_check_76_to_variable;

// 拆分后校验节点76传递给变量节点14的值以及对变量节点14传递过来的值
wire [5:0] value_check_76_to_variable_14;
wire enable_check_76_to_variable_14;
wire [5:0] value_variable_14_to_check_76;
wire enable_variable_14_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_14 = value_check_76_to_variable[5:0];
assign enable_check_76_to_variable_14 = enable_check_76_to_variable[0];
// 对变量节点14传递过来的值进行组合
assign value_variable_to_check_76[5:0] = value_variable_14_to_check_76;
assign enable_variable_to_check_76[0] = enable_variable_14_to_check_76;

// 拆分后校验节点76传递给变量节点63的值以及对变量节点63传递过来的值
wire [5:0] value_check_76_to_variable_63;
wire enable_check_76_to_variable_63;
wire [5:0] value_variable_63_to_check_76;
wire enable_variable_63_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_63 = value_check_76_to_variable[11:6];
assign enable_check_76_to_variable_63 = enable_check_76_to_variable[1];
// 对变量节点63传递过来的值进行组合
assign value_variable_to_check_76[11:6] = value_variable_63_to_check_76;
assign enable_variable_to_check_76[1] = enable_variable_63_to_check_76;

// 拆分后校验节点76传递给变量节点105的值以及对变量节点105传递过来的值
wire [5:0] value_check_76_to_variable_105;
wire enable_check_76_to_variable_105;
wire [5:0] value_variable_105_to_check_76;
wire enable_variable_105_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_105 = value_check_76_to_variable[17:12];
assign enable_check_76_to_variable_105 = enable_check_76_to_variable[2];
// 对变量节点105传递过来的值进行组合
assign value_variable_to_check_76[17:12] = value_variable_105_to_check_76;
assign enable_variable_to_check_76[2] = enable_variable_105_to_check_76;

// 拆分后校验节点76传递给变量节点131的值以及对变量节点131传递过来的值
wire [5:0] value_check_76_to_variable_131;
wire enable_check_76_to_variable_131;
wire [5:0] value_variable_131_to_check_76;
wire enable_variable_131_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_131 = value_check_76_to_variable[23:18];
assign enable_check_76_to_variable_131 = enable_check_76_to_variable[3];
// 对变量节点131传递过来的值进行组合
assign value_variable_to_check_76[23:18] = value_variable_131_to_check_76;
assign enable_variable_to_check_76[3] = enable_variable_131_to_check_76;

// 拆分后校验节点76传递给变量节点194的值以及对变量节点194传递过来的值
wire [5:0] value_check_76_to_variable_194;
wire enable_check_76_to_variable_194;
wire [5:0] value_variable_194_to_check_76;
wire enable_variable_194_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_194 = value_check_76_to_variable[29:24];
assign enable_check_76_to_variable_194 = enable_check_76_to_variable[4];
// 对变量节点194传递过来的值进行组合
assign value_variable_to_check_76[29:24] = value_variable_194_to_check_76;
assign enable_variable_to_check_76[4] = enable_variable_194_to_check_76;

// 拆分后校验节点76传递给变量节点253的值以及对变量节点253传递过来的值
wire [5:0] value_check_76_to_variable_253;
wire enable_check_76_to_variable_253;
wire [5:0] value_variable_253_to_check_76;
wire enable_variable_253_to_check_76;
// 对校验节点76的输出值进行拆分
assign value_check_76_to_variable_253 = value_check_76_to_variable[35:30];
assign enable_check_76_to_variable_253 = enable_check_76_to_variable[5];
// 对变量节点253传递过来的值进行组合
assign value_variable_to_check_76[35:30] = value_variable_253_to_check_76;
assign enable_variable_to_check_76[5] = enable_variable_253_to_check_76;


// 校验节点77的接口
wire [35:0] value_variable_to_check_77;
wire [35:0] value_check_77_to_variable;
wire [5:0] enable_variable_to_check_77;
wire [5:0] enable_check_77_to_variable;

// 拆分后校验节点77传递给变量节点37的值以及对变量节点37传递过来的值
wire [5:0] value_check_77_to_variable_37;
wire enable_check_77_to_variable_37;
wire [5:0] value_variable_37_to_check_77;
wire enable_variable_37_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_37 = value_check_77_to_variable[5:0];
assign enable_check_77_to_variable_37 = enable_check_77_to_variable[0];
// 对变量节点37传递过来的值进行组合
assign value_variable_to_check_77[5:0] = value_variable_37_to_check_77;
assign enable_variable_to_check_77[0] = enable_variable_37_to_check_77;

// 拆分后校验节点77传递给变量节点50的值以及对变量节点50传递过来的值
wire [5:0] value_check_77_to_variable_50;
wire enable_check_77_to_variable_50;
wire [5:0] value_variable_50_to_check_77;
wire enable_variable_50_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_50 = value_check_77_to_variable[11:6];
assign enable_check_77_to_variable_50 = enable_check_77_to_variable[1];
// 对变量节点50传递过来的值进行组合
assign value_variable_to_check_77[11:6] = value_variable_50_to_check_77;
assign enable_variable_to_check_77[1] = enable_variable_50_to_check_77;

// 拆分后校验节点77传递给变量节点107的值以及对变量节点107传递过来的值
wire [5:0] value_check_77_to_variable_107;
wire enable_check_77_to_variable_107;
wire [5:0] value_variable_107_to_check_77;
wire enable_variable_107_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_107 = value_check_77_to_variable[17:12];
assign enable_check_77_to_variable_107 = enable_check_77_to_variable[2];
// 对变量节点107传递过来的值进行组合
assign value_variable_to_check_77[17:12] = value_variable_107_to_check_77;
assign enable_variable_to_check_77[2] = enable_variable_107_to_check_77;

// 拆分后校验节点77传递给变量节点140的值以及对变量节点140传递过来的值
wire [5:0] value_check_77_to_variable_140;
wire enable_check_77_to_variable_140;
wire [5:0] value_variable_140_to_check_77;
wire enable_variable_140_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_140 = value_check_77_to_variable[23:18];
assign enable_check_77_to_variable_140 = enable_check_77_to_variable[3];
// 对变量节点140传递过来的值进行组合
assign value_variable_to_check_77[23:18] = value_variable_140_to_check_77;
assign enable_variable_to_check_77[3] = enable_variable_140_to_check_77;

// 拆分后校验节点77传递给变量节点205的值以及对变量节点205传递过来的值
wire [5:0] value_check_77_to_variable_205;
wire enable_check_77_to_variable_205;
wire [5:0] value_variable_205_to_check_77;
wire enable_variable_205_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_205 = value_check_77_to_variable[29:24];
assign enable_check_77_to_variable_205 = enable_check_77_to_variable[4];
// 对变量节点205传递过来的值进行组合
assign value_variable_to_check_77[29:24] = value_variable_205_to_check_77;
assign enable_variable_to_check_77[4] = enable_variable_205_to_check_77;

// 拆分后校验节点77传递给变量节点245的值以及对变量节点245传递过来的值
wire [5:0] value_check_77_to_variable_245;
wire enable_check_77_to_variable_245;
wire [5:0] value_variable_245_to_check_77;
wire enable_variable_245_to_check_77;
// 对校验节点77的输出值进行拆分
assign value_check_77_to_variable_245 = value_check_77_to_variable[35:30];
assign enable_check_77_to_variable_245 = enable_check_77_to_variable[5];
// 对变量节点245传递过来的值进行组合
assign value_variable_to_check_77[35:30] = value_variable_245_to_check_77;
assign enable_variable_to_check_77[5] = enable_variable_245_to_check_77;


// 校验节点78的接口
wire [35:0] value_variable_to_check_78;
wire [35:0] value_check_78_to_variable;
wire [5:0] enable_variable_to_check_78;
wire [5:0] enable_check_78_to_variable;

// 拆分后校验节点78传递给变量节点33的值以及对变量节点33传递过来的值
wire [5:0] value_check_78_to_variable_33;
wire enable_check_78_to_variable_33;
wire [5:0] value_variable_33_to_check_78;
wire enable_variable_33_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_33 = value_check_78_to_variable[5:0];
assign enable_check_78_to_variable_33 = enable_check_78_to_variable[0];
// 对变量节点33传递过来的值进行组合
assign value_variable_to_check_78[5:0] = value_variable_33_to_check_78;
assign enable_variable_to_check_78[0] = enable_variable_33_to_check_78;

// 拆分后校验节点78传递给变量节点49的值以及对变量节点49传递过来的值
wire [5:0] value_check_78_to_variable_49;
wire enable_check_78_to_variable_49;
wire [5:0] value_variable_49_to_check_78;
wire enable_variable_49_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_49 = value_check_78_to_variable[11:6];
assign enable_check_78_to_variable_49 = enable_check_78_to_variable[1];
// 对变量节点49传递过来的值进行组合
assign value_variable_to_check_78[11:6] = value_variable_49_to_check_78;
assign enable_variable_to_check_78[1] = enable_variable_49_to_check_78;

// 拆分后校验节点78传递给变量节点97的值以及对变量节点97传递过来的值
wire [5:0] value_check_78_to_variable_97;
wire enable_check_78_to_variable_97;
wire [5:0] value_variable_97_to_check_78;
wire enable_variable_97_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_97 = value_check_78_to_variable[17:12];
assign enable_check_78_to_variable_97 = enable_check_78_to_variable[2];
// 对变量节点97传递过来的值进行组合
assign value_variable_to_check_78[17:12] = value_variable_97_to_check_78;
assign enable_variable_to_check_78[2] = enable_variable_97_to_check_78;

// 拆分后校验节点78传递给变量节点109的值以及对变量节点109传递过来的值
wire [5:0] value_check_78_to_variable_109;
wire enable_check_78_to_variable_109;
wire [5:0] value_variable_109_to_check_78;
wire enable_variable_109_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_109 = value_check_78_to_variable[23:18];
assign enable_check_78_to_variable_109 = enable_check_78_to_variable[3];
// 对变量节点109传递过来的值进行组合
assign value_variable_to_check_78[23:18] = value_variable_109_to_check_78;
assign enable_variable_to_check_78[3] = enable_variable_109_to_check_78;

// 拆分后校验节点78传递给变量节点186的值以及对变量节点186传递过来的值
wire [5:0] value_check_78_to_variable_186;
wire enable_check_78_to_variable_186;
wire [5:0] value_variable_186_to_check_78;
wire enable_variable_186_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_186 = value_check_78_to_variable[29:24];
assign enable_check_78_to_variable_186 = enable_check_78_to_variable[4];
// 对变量节点186传递过来的值进行组合
assign value_variable_to_check_78[29:24] = value_variable_186_to_check_78;
assign enable_variable_to_check_78[4] = enable_variable_186_to_check_78;

// 拆分后校验节点78传递给变量节点218的值以及对变量节点218传递过来的值
wire [5:0] value_check_78_to_variable_218;
wire enable_check_78_to_variable_218;
wire [5:0] value_variable_218_to_check_78;
wire enable_variable_218_to_check_78;
// 对校验节点78的输出值进行拆分
assign value_check_78_to_variable_218 = value_check_78_to_variable[35:30];
assign enable_check_78_to_variable_218 = enable_check_78_to_variable[5];
// 对变量节点218传递过来的值进行组合
assign value_variable_to_check_78[35:30] = value_variable_218_to_check_78;
assign enable_variable_to_check_78[5] = enable_variable_218_to_check_78;


// 校验节点79的接口
wire [35:0] value_variable_to_check_79;
wire [35:0] value_check_79_to_variable;
wire [5:0] enable_variable_to_check_79;
wire [5:0] enable_check_79_to_variable;

// 拆分后校验节点79传递给变量节点39的值以及对变量节点39传递过来的值
wire [5:0] value_check_79_to_variable_39;
wire enable_check_79_to_variable_39;
wire [5:0] value_variable_39_to_check_79;
wire enable_variable_39_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_39 = value_check_79_to_variable[5:0];
assign enable_check_79_to_variable_39 = enable_check_79_to_variable[0];
// 对变量节点39传递过来的值进行组合
assign value_variable_to_check_79[5:0] = value_variable_39_to_check_79;
assign enable_variable_to_check_79[0] = enable_variable_39_to_check_79;

// 拆分后校验节点79传递给变量节点78的值以及对变量节点78传递过来的值
wire [5:0] value_check_79_to_variable_78;
wire enable_check_79_to_variable_78;
wire [5:0] value_variable_78_to_check_79;
wire enable_variable_78_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_78 = value_check_79_to_variable[11:6];
assign enable_check_79_to_variable_78 = enable_check_79_to_variable[1];
// 对变量节点78传递过来的值进行组合
assign value_variable_to_check_79[11:6] = value_variable_78_to_check_79;
assign enable_variable_to_check_79[1] = enable_variable_78_to_check_79;

// 拆分后校验节点79传递给变量节点111的值以及对变量节点111传递过来的值
wire [5:0] value_check_79_to_variable_111;
wire enable_check_79_to_variable_111;
wire [5:0] value_variable_111_to_check_79;
wire enable_variable_111_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_111 = value_check_79_to_variable[17:12];
assign enable_check_79_to_variable_111 = enable_check_79_to_variable[2];
// 对变量节点111传递过来的值进行组合
assign value_variable_to_check_79[17:12] = value_variable_111_to_check_79;
assign enable_variable_to_check_79[2] = enable_variable_111_to_check_79;

// 拆分后校验节点79传递给变量节点163的值以及对变量节点163传递过来的值
wire [5:0] value_check_79_to_variable_163;
wire enable_check_79_to_variable_163;
wire [5:0] value_variable_163_to_check_79;
wire enable_variable_163_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_163 = value_check_79_to_variable[23:18];
assign enable_check_79_to_variable_163 = enable_check_79_to_variable[3];
// 对变量节点163传递过来的值进行组合
assign value_variable_to_check_79[23:18] = value_variable_163_to_check_79;
assign enable_variable_to_check_79[3] = enable_variable_163_to_check_79;

// 拆分后校验节点79传递给变量节点210的值以及对变量节点210传递过来的值
wire [5:0] value_check_79_to_variable_210;
wire enable_check_79_to_variable_210;
wire [5:0] value_variable_210_to_check_79;
wire enable_variable_210_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_210 = value_check_79_to_variable[29:24];
assign enable_check_79_to_variable_210 = enable_check_79_to_variable[4];
// 对变量节点210传递过来的值进行组合
assign value_variable_to_check_79[29:24] = value_variable_210_to_check_79;
assign enable_variable_to_check_79[4] = enable_variable_210_to_check_79;

// 拆分后校验节点79传递给变量节点242的值以及对变量节点242传递过来的值
wire [5:0] value_check_79_to_variable_242;
wire enable_check_79_to_variable_242;
wire [5:0] value_variable_242_to_check_79;
wire enable_variable_242_to_check_79;
// 对校验节点79的输出值进行拆分
assign value_check_79_to_variable_242 = value_check_79_to_variable[35:30];
assign enable_check_79_to_variable_242 = enable_check_79_to_variable[5];
// 对变量节点242传递过来的值进行组合
assign value_variable_to_check_79[35:30] = value_variable_242_to_check_79;
assign enable_variable_to_check_79[5] = enable_variable_242_to_check_79;


// 校验节点80的接口
wire [35:0] value_variable_to_check_80;
wire [35:0] value_check_80_to_variable;
wire [5:0] enable_variable_to_check_80;
wire [5:0] enable_check_80_to_variable;

// 拆分后校验节点80传递给变量节点35的值以及对变量节点35传递过来的值
wire [5:0] value_check_80_to_variable_35;
wire enable_check_80_to_variable_35;
wire [5:0] value_variable_35_to_check_80;
wire enable_variable_35_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_35 = value_check_80_to_variable[5:0];
assign enable_check_80_to_variable_35 = enable_check_80_to_variable[0];
// 对变量节点35传递过来的值进行组合
assign value_variable_to_check_80[5:0] = value_variable_35_to_check_80;
assign enable_variable_to_check_80[0] = enable_variable_35_to_check_80;

// 拆分后校验节点80传递给变量节点43的值以及对变量节点43传递过来的值
wire [5:0] value_check_80_to_variable_43;
wire enable_check_80_to_variable_43;
wire [5:0] value_variable_43_to_check_80;
wire enable_variable_43_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_43 = value_check_80_to_variable[11:6];
assign enable_check_80_to_variable_43 = enable_check_80_to_variable[1];
// 对变量节点43传递过来的值进行组合
assign value_variable_to_check_80[11:6] = value_variable_43_to_check_80;
assign enable_variable_to_check_80[1] = enable_variable_43_to_check_80;

// 拆分后校验节点80传递给变量节点122的值以及对变量节点122传递过来的值
wire [5:0] value_check_80_to_variable_122;
wire enable_check_80_to_variable_122;
wire [5:0] value_variable_122_to_check_80;
wire enable_variable_122_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_122 = value_check_80_to_variable[17:12];
assign enable_check_80_to_variable_122 = enable_check_80_to_variable[2];
// 对变量节点122传递过来的值进行组合
assign value_variable_to_check_80[17:12] = value_variable_122_to_check_80;
assign enable_variable_to_check_80[2] = enable_variable_122_to_check_80;

// 拆分后校验节点80传递给变量节点155的值以及对变量节点155传递过来的值
wire [5:0] value_check_80_to_variable_155;
wire enable_check_80_to_variable_155;
wire [5:0] value_variable_155_to_check_80;
wire enable_variable_155_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_155 = value_check_80_to_variable[23:18];
assign enable_check_80_to_variable_155 = enable_check_80_to_variable[3];
// 对变量节点155传递过来的值进行组合
assign value_variable_to_check_80[23:18] = value_variable_155_to_check_80;
assign enable_variable_to_check_80[3] = enable_variable_155_to_check_80;

// 拆分后校验节点80传递给变量节点201的值以及对变量节点201传递过来的值
wire [5:0] value_check_80_to_variable_201;
wire enable_check_80_to_variable_201;
wire [5:0] value_variable_201_to_check_80;
wire enable_variable_201_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_201 = value_check_80_to_variable[29:24];
assign enable_check_80_to_variable_201 = enable_check_80_to_variable[4];
// 对变量节点201传递过来的值进行组合
assign value_variable_to_check_80[29:24] = value_variable_201_to_check_80;
assign enable_variable_to_check_80[4] = enable_variable_201_to_check_80;

// 拆分后校验节点80传递给变量节点254的值以及对变量节点254传递过来的值
wire [5:0] value_check_80_to_variable_254;
wire enable_check_80_to_variable_254;
wire [5:0] value_variable_254_to_check_80;
wire enable_variable_254_to_check_80;
// 对校验节点80的输出值进行拆分
assign value_check_80_to_variable_254 = value_check_80_to_variable[35:30];
assign enable_check_80_to_variable_254 = enable_check_80_to_variable[5];
// 对变量节点254传递过来的值进行组合
assign value_variable_to_check_80[35:30] = value_variable_254_to_check_80;
assign enable_variable_to_check_80[5] = enable_variable_254_to_check_80;


// 校验节点81的接口
wire [35:0] value_variable_to_check_81;
wire [35:0] value_check_81_to_variable;
wire [5:0] enable_variable_to_check_81;
wire [5:0] enable_check_81_to_variable;

// 拆分后校验节点81传递给变量节点13的值以及对变量节点13传递过来的值
wire [5:0] value_check_81_to_variable_13;
wire enable_check_81_to_variable_13;
wire [5:0] value_variable_13_to_check_81;
wire enable_variable_13_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_13 = value_check_81_to_variable[5:0];
assign enable_check_81_to_variable_13 = enable_check_81_to_variable[0];
// 对变量节点13传递过来的值进行组合
assign value_variable_to_check_81[5:0] = value_variable_13_to_check_81;
assign enable_variable_to_check_81[0] = enable_variable_13_to_check_81;

// 拆分后校验节点81传递给变量节点76的值以及对变量节点76传递过来的值
wire [5:0] value_check_81_to_variable_76;
wire enable_check_81_to_variable_76;
wire [5:0] value_variable_76_to_check_81;
wire enable_variable_76_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_76 = value_check_81_to_variable[11:6];
assign enable_check_81_to_variable_76 = enable_check_81_to_variable[1];
// 对变量节点76传递过来的值进行组合
assign value_variable_to_check_81[11:6] = value_variable_76_to_check_81;
assign enable_variable_to_check_81[1] = enable_variable_76_to_check_81;

// 拆分后校验节点81传递给变量节点124的值以及对变量节点124传递过来的值
wire [5:0] value_check_81_to_variable_124;
wire enable_check_81_to_variable_124;
wire [5:0] value_variable_124_to_check_81;
wire enable_variable_124_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_124 = value_check_81_to_variable[17:12];
assign enable_check_81_to_variable_124 = enable_check_81_to_variable[2];
// 对变量节点124传递过来的值进行组合
assign value_variable_to_check_81[17:12] = value_variable_124_to_check_81;
assign enable_variable_to_check_81[2] = enable_variable_124_to_check_81;

// 拆分后校验节点81传递给变量节点148的值以及对变量节点148传递过来的值
wire [5:0] value_check_81_to_variable_148;
wire enable_check_81_to_variable_148;
wire [5:0] value_variable_148_to_check_81;
wire enable_variable_148_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_148 = value_check_81_to_variable[23:18];
assign enable_check_81_to_variable_148 = enable_check_81_to_variable[3];
// 对变量节点148传递过来的值进行组合
assign value_variable_to_check_81[23:18] = value_variable_148_to_check_81;
assign enable_variable_to_check_81[3] = enable_variable_148_to_check_81;

// 拆分后校验节点81传递给变量节点201的值以及对变量节点201传递过来的值
wire [5:0] value_check_81_to_variable_201;
wire enable_check_81_to_variable_201;
wire [5:0] value_variable_201_to_check_81;
wire enable_variable_201_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_201 = value_check_81_to_variable[29:24];
assign enable_check_81_to_variable_201 = enable_check_81_to_variable[4];
// 对变量节点201传递过来的值进行组合
assign value_variable_to_check_81[29:24] = value_variable_201_to_check_81;
assign enable_variable_to_check_81[4] = enable_variable_201_to_check_81;

// 拆分后校验节点81传递给变量节点234的值以及对变量节点234传递过来的值
wire [5:0] value_check_81_to_variable_234;
wire enable_check_81_to_variable_234;
wire [5:0] value_variable_234_to_check_81;
wire enable_variable_234_to_check_81;
// 对校验节点81的输出值进行拆分
assign value_check_81_to_variable_234 = value_check_81_to_variable[35:30];
assign enable_check_81_to_variable_234 = enable_check_81_to_variable[5];
// 对变量节点234传递过来的值进行组合
assign value_variable_to_check_81[35:30] = value_variable_234_to_check_81;
assign enable_variable_to_check_81[5] = enable_variable_234_to_check_81;


// 校验节点82的接口
wire [35:0] value_variable_to_check_82;
wire [35:0] value_check_82_to_variable;
wire [5:0] enable_variable_to_check_82;
wire [5:0] enable_check_82_to_variable;

// 拆分后校验节点82传递给变量节点41的值以及对变量节点41传递过来的值
wire [5:0] value_check_82_to_variable_41;
wire enable_check_82_to_variable_41;
wire [5:0] value_variable_41_to_check_82;
wire enable_variable_41_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_41 = value_check_82_to_variable[5:0];
assign enable_check_82_to_variable_41 = enable_check_82_to_variable[0];
// 对变量节点41传递过来的值进行组合
assign value_variable_to_check_82[5:0] = value_variable_41_to_check_82;
assign enable_variable_to_check_82[0] = enable_variable_41_to_check_82;

// 拆分后校验节点82传递给变量节点82的值以及对变量节点82传递过来的值
wire [5:0] value_check_82_to_variable_82;
wire enable_check_82_to_variable_82;
wire [5:0] value_variable_82_to_check_82;
wire enable_variable_82_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_82 = value_check_82_to_variable[11:6];
assign enable_check_82_to_variable_82 = enable_check_82_to_variable[1];
// 对变量节点82传递过来的值进行组合
assign value_variable_to_check_82[11:6] = value_variable_82_to_check_82;
assign enable_variable_to_check_82[1] = enable_variable_82_to_check_82;

// 拆分后校验节点82传递给变量节点125的值以及对变量节点125传递过来的值
wire [5:0] value_check_82_to_variable_125;
wire enable_check_82_to_variable_125;
wire [5:0] value_variable_125_to_check_82;
wire enable_variable_125_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_125 = value_check_82_to_variable[17:12];
assign enable_check_82_to_variable_125 = enable_check_82_to_variable[2];
// 对变量节点125传递过来的值进行组合
assign value_variable_to_check_82[17:12] = value_variable_125_to_check_82;
assign enable_variable_to_check_82[2] = enable_variable_125_to_check_82;

// 拆分后校验节点82传递给变量节点164的值以及对变量节点164传递过来的值
wire [5:0] value_check_82_to_variable_164;
wire enable_check_82_to_variable_164;
wire [5:0] value_variable_164_to_check_82;
wire enable_variable_164_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_164 = value_check_82_to_variable[23:18];
assign enable_check_82_to_variable_164 = enable_check_82_to_variable[3];
// 对变量节点164传递过来的值进行组合
assign value_variable_to_check_82[23:18] = value_variable_164_to_check_82;
assign enable_variable_to_check_82[3] = enable_variable_164_to_check_82;

// 拆分后校验节点82传递给变量节点176的值以及对变量节点176传递过来的值
wire [5:0] value_check_82_to_variable_176;
wire enable_check_82_to_variable_176;
wire [5:0] value_variable_176_to_check_82;
wire enable_variable_176_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_176 = value_check_82_to_variable[29:24];
assign enable_check_82_to_variable_176 = enable_check_82_to_variable[4];
// 对变量节点176传递过来的值进行组合
assign value_variable_to_check_82[29:24] = value_variable_176_to_check_82;
assign enable_variable_to_check_82[4] = enable_variable_176_to_check_82;

// 拆分后校验节点82传递给变量节点252的值以及对变量节点252传递过来的值
wire [5:0] value_check_82_to_variable_252;
wire enable_check_82_to_variable_252;
wire [5:0] value_variable_252_to_check_82;
wire enable_variable_252_to_check_82;
// 对校验节点82的输出值进行拆分
assign value_check_82_to_variable_252 = value_check_82_to_variable[35:30];
assign enable_check_82_to_variable_252 = enable_check_82_to_variable[5];
// 对变量节点252传递过来的值进行组合
assign value_variable_to_check_82[35:30] = value_variable_252_to_check_82;
assign enable_variable_to_check_82[5] = enable_variable_252_to_check_82;


// 校验节点83的接口
wire [35:0] value_variable_to_check_83;
wire [35:0] value_check_83_to_variable;
wire [5:0] enable_variable_to_check_83;
wire [5:0] enable_check_83_to_variable;

// 拆分后校验节点83传递给变量节点29的值以及对变量节点29传递过来的值
wire [5:0] value_check_83_to_variable_29;
wire enable_check_83_to_variable_29;
wire [5:0] value_variable_29_to_check_83;
wire enable_variable_29_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_29 = value_check_83_to_variable[5:0];
assign enable_check_83_to_variable_29 = enable_check_83_to_variable[0];
// 对变量节点29传递过来的值进行组合
assign value_variable_to_check_83[5:0] = value_variable_29_to_check_83;
assign enable_variable_to_check_83[0] = enable_variable_29_to_check_83;

// 拆分后校验节点83传递给变量节点55的值以及对变量节点55传递过来的值
wire [5:0] value_check_83_to_variable_55;
wire enable_check_83_to_variable_55;
wire [5:0] value_variable_55_to_check_83;
wire enable_variable_55_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_55 = value_check_83_to_variable[11:6];
assign enable_check_83_to_variable_55 = enable_check_83_to_variable[1];
// 对变量节点55传递过来的值进行组合
assign value_variable_to_check_83[11:6] = value_variable_55_to_check_83;
assign enable_variable_to_check_83[1] = enable_variable_55_to_check_83;

// 拆分后校验节点83传递给变量节点126的值以及对变量节点126传递过来的值
wire [5:0] value_check_83_to_variable_126;
wire enable_check_83_to_variable_126;
wire [5:0] value_variable_126_to_check_83;
wire enable_variable_126_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_126 = value_check_83_to_variable[17:12];
assign enable_check_83_to_variable_126 = enable_check_83_to_variable[2];
// 对变量节点126传递过来的值进行组合
assign value_variable_to_check_83[17:12] = value_variable_126_to_check_83;
assign enable_variable_to_check_83[2] = enable_variable_126_to_check_83;

// 拆分后校验节点83传递给变量节点140的值以及对变量节点140传递过来的值
wire [5:0] value_check_83_to_variable_140;
wire enable_check_83_to_variable_140;
wire [5:0] value_variable_140_to_check_83;
wire enable_variable_140_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_140 = value_check_83_to_variable[23:18];
assign enable_check_83_to_variable_140 = enable_check_83_to_variable[3];
// 对变量节点140传递过来的值进行组合
assign value_variable_to_check_83[23:18] = value_variable_140_to_check_83;
assign enable_variable_to_check_83[3] = enable_variable_140_to_check_83;

// 拆分后校验节点83传递给变量节点203的值以及对变量节点203传递过来的值
wire [5:0] value_check_83_to_variable_203;
wire enable_check_83_to_variable_203;
wire [5:0] value_variable_203_to_check_83;
wire enable_variable_203_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_203 = value_check_83_to_variable[29:24];
assign enable_check_83_to_variable_203 = enable_check_83_to_variable[4];
// 对变量节点203传递过来的值进行组合
assign value_variable_to_check_83[29:24] = value_variable_203_to_check_83;
assign enable_variable_to_check_83[4] = enable_variable_203_to_check_83;

// 拆分后校验节点83传递给变量节点220的值以及对变量节点220传递过来的值
wire [5:0] value_check_83_to_variable_220;
wire enable_check_83_to_variable_220;
wire [5:0] value_variable_220_to_check_83;
wire enable_variable_220_to_check_83;
// 对校验节点83的输出值进行拆分
assign value_check_83_to_variable_220 = value_check_83_to_variable[35:30];
assign enable_check_83_to_variable_220 = enable_check_83_to_variable[5];
// 对变量节点220传递过来的值进行组合
assign value_variable_to_check_83[35:30] = value_variable_220_to_check_83;
assign enable_variable_to_check_83[5] = enable_variable_220_to_check_83;


// 校验节点84的接口
wire [35:0] value_variable_to_check_84;
wire [35:0] value_check_84_to_variable;
wire [5:0] enable_variable_to_check_84;
wire [5:0] enable_check_84_to_variable;

// 拆分后校验节点84传递给变量节点28的值以及对变量节点28传递过来的值
wire [5:0] value_check_84_to_variable_28;
wire enable_check_84_to_variable_28;
wire [5:0] value_variable_28_to_check_84;
wire enable_variable_28_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_28 = value_check_84_to_variable[5:0];
assign enable_check_84_to_variable_28 = enable_check_84_to_variable[0];
// 对变量节点28传递过来的值进行组合
assign value_variable_to_check_84[5:0] = value_variable_28_to_check_84;
assign enable_variable_to_check_84[0] = enable_variable_28_to_check_84;

// 拆分后校验节点84传递给变量节点68的值以及对变量节点68传递过来的值
wire [5:0] value_check_84_to_variable_68;
wire enable_check_84_to_variable_68;
wire [5:0] value_variable_68_to_check_84;
wire enable_variable_68_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_68 = value_check_84_to_variable[11:6];
assign enable_check_84_to_variable_68 = enable_check_84_to_variable[1];
// 对变量节点68传递过来的值进行组合
assign value_variable_to_check_84[11:6] = value_variable_68_to_check_84;
assign enable_variable_to_check_84[1] = enable_variable_68_to_check_84;

// 拆分后校验节点84传递给变量节点116的值以及对变量节点116传递过来的值
wire [5:0] value_check_84_to_variable_116;
wire enable_check_84_to_variable_116;
wire [5:0] value_variable_116_to_check_84;
wire enable_variable_116_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_116 = value_check_84_to_variable[17:12];
assign enable_check_84_to_variable_116 = enable_check_84_to_variable[2];
// 对变量节点116传递过来的值进行组合
assign value_variable_to_check_84[17:12] = value_variable_116_to_check_84;
assign enable_variable_to_check_84[2] = enable_variable_116_to_check_84;

// 拆分后校验节点84传递给变量节点159的值以及对变量节点159传递过来的值
wire [5:0] value_check_84_to_variable_159;
wire enable_check_84_to_variable_159;
wire [5:0] value_variable_159_to_check_84;
wire enable_variable_159_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_159 = value_check_84_to_variable[23:18];
assign enable_check_84_to_variable_159 = enable_check_84_to_variable[3];
// 对变量节点159传递过来的值进行组合
assign value_variable_to_check_84[23:18] = value_variable_159_to_check_84;
assign enable_variable_to_check_84[3] = enable_variable_159_to_check_84;

// 拆分后校验节点84传递给变量节点209的值以及对变量节点209传递过来的值
wire [5:0] value_check_84_to_variable_209;
wire enable_check_84_to_variable_209;
wire [5:0] value_variable_209_to_check_84;
wire enable_variable_209_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_209 = value_check_84_to_variable[29:24];
assign enable_check_84_to_variable_209 = enable_check_84_to_variable[4];
// 对变量节点209传递过来的值进行组合
assign value_variable_to_check_84[29:24] = value_variable_209_to_check_84;
assign enable_variable_to_check_84[4] = enable_variable_209_to_check_84;

// 拆分后校验节点84传递给变量节点243的值以及对变量节点243传递过来的值
wire [5:0] value_check_84_to_variable_243;
wire enable_check_84_to_variable_243;
wire [5:0] value_variable_243_to_check_84;
wire enable_variable_243_to_check_84;
// 对校验节点84的输出值进行拆分
assign value_check_84_to_variable_243 = value_check_84_to_variable[35:30];
assign enable_check_84_to_variable_243 = enable_check_84_to_variable[5];
// 对变量节点243传递过来的值进行组合
assign value_variable_to_check_84[35:30] = value_variable_243_to_check_84;
assign enable_variable_to_check_84[5] = enable_variable_243_to_check_84;


// 校验节点85的接口
wire [35:0] value_variable_to_check_85;
wire [35:0] value_check_85_to_variable;
wire [5:0] enable_variable_to_check_85;
wire [5:0] enable_check_85_to_variable;

// 拆分后校验节点85传递给变量节点25的值以及对变量节点25传递过来的值
wire [5:0] value_check_85_to_variable_25;
wire enable_check_85_to_variable_25;
wire [5:0] value_variable_25_to_check_85;
wire enable_variable_25_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_25 = value_check_85_to_variable[5:0];
assign enable_check_85_to_variable_25 = enable_check_85_to_variable[0];
// 对变量节点25传递过来的值进行组合
assign value_variable_to_check_85[5:0] = value_variable_25_to_check_85;
assign enable_variable_to_check_85[0] = enable_variable_25_to_check_85;

// 拆分后校验节点85传递给变量节点77的值以及对变量节点77传递过来的值
wire [5:0] value_check_85_to_variable_77;
wire enable_check_85_to_variable_77;
wire [5:0] value_variable_77_to_check_85;
wire enable_variable_77_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_77 = value_check_85_to_variable[11:6];
assign enable_check_85_to_variable_77 = enable_check_85_to_variable[1];
// 对变量节点77传递过来的值进行组合
assign value_variable_to_check_85[11:6] = value_variable_77_to_check_85;
assign enable_variable_to_check_85[1] = enable_variable_77_to_check_85;

// 拆分后校验节点85传递给变量节点127的值以及对变量节点127传递过来的值
wire [5:0] value_check_85_to_variable_127;
wire enable_check_85_to_variable_127;
wire [5:0] value_variable_127_to_check_85;
wire enable_variable_127_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_127 = value_check_85_to_variable[17:12];
assign enable_check_85_to_variable_127 = enable_check_85_to_variable[2];
// 对变量节点127传递过来的值进行组合
assign value_variable_to_check_85[17:12] = value_variable_127_to_check_85;
assign enable_variable_to_check_85[2] = enable_variable_127_to_check_85;

// 拆分后校验节点85传递给变量节点129的值以及对变量节点129传递过来的值
wire [5:0] value_check_85_to_variable_129;
wire enable_check_85_to_variable_129;
wire [5:0] value_variable_129_to_check_85;
wire enable_variable_129_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_129 = value_check_85_to_variable[23:18];
assign enable_check_85_to_variable_129 = enable_check_85_to_variable[3];
// 对变量节点129传递过来的值进行组合
assign value_variable_to_check_85[23:18] = value_variable_129_to_check_85;
assign enable_variable_to_check_85[3] = enable_variable_129_to_check_85;

// 拆分后校验节点85传递给变量节点183的值以及对变量节点183传递过来的值
wire [5:0] value_check_85_to_variable_183;
wire enable_check_85_to_variable_183;
wire [5:0] value_variable_183_to_check_85;
wire enable_variable_183_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_183 = value_check_85_to_variable[29:24];
assign enable_check_85_to_variable_183 = enable_check_85_to_variable[4];
// 对变量节点183传递过来的值进行组合
assign value_variable_to_check_85[29:24] = value_variable_183_to_check_85;
assign enable_variable_to_check_85[4] = enable_variable_183_to_check_85;

// 拆分后校验节点85传递给变量节点250的值以及对变量节点250传递过来的值
wire [5:0] value_check_85_to_variable_250;
wire enable_check_85_to_variable_250;
wire [5:0] value_variable_250_to_check_85;
wire enable_variable_250_to_check_85;
// 对校验节点85的输出值进行拆分
assign value_check_85_to_variable_250 = value_check_85_to_variable[35:30];
assign enable_check_85_to_variable_250 = enable_check_85_to_variable[5];
// 对变量节点250传递过来的值进行组合
assign value_variable_to_check_85[35:30] = value_variable_250_to_check_85;
assign enable_variable_to_check_85[5] = enable_variable_250_to_check_85;


// 校验节点86的接口
wire [35:0] value_variable_to_check_86;
wire [35:0] value_check_86_to_variable;
wire [5:0] enable_variable_to_check_86;
wire [5:0] enable_check_86_to_variable;

// 拆分后校验节点86传递给变量节点35的值以及对变量节点35传递过来的值
wire [5:0] value_check_86_to_variable_35;
wire enable_check_86_to_variable_35;
wire [5:0] value_variable_35_to_check_86;
wire enable_variable_35_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_35 = value_check_86_to_variable[5:0];
assign enable_check_86_to_variable_35 = enable_check_86_to_variable[0];
// 对变量节点35传递过来的值进行组合
assign value_variable_to_check_86[5:0] = value_variable_35_to_check_86;
assign enable_variable_to_check_86[0] = enable_variable_35_to_check_86;

// 拆分后校验节点86传递给变量节点47的值以及对变量节点47传递过来的值
wire [5:0] value_check_86_to_variable_47;
wire enable_check_86_to_variable_47;
wire [5:0] value_variable_47_to_check_86;
wire enable_variable_47_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_47 = value_check_86_to_variable[11:6];
assign enable_check_86_to_variable_47 = enable_check_86_to_variable[1];
// 对变量节点47传递过来的值进行组合
assign value_variable_to_check_86[11:6] = value_variable_47_to_check_86;
assign enable_variable_to_check_86[1] = enable_variable_47_to_check_86;

// 拆分后校验节点86传递给变量节点128的值以及对变量节点128传递过来的值
wire [5:0] value_check_86_to_variable_128;
wire enable_check_86_to_variable_128;
wire [5:0] value_variable_128_to_check_86;
wire enable_variable_128_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_128 = value_check_86_to_variable[17:12];
assign enable_check_86_to_variable_128 = enable_check_86_to_variable[2];
// 对变量节点128传递过来的值进行组合
assign value_variable_to_check_86[17:12] = value_variable_128_to_check_86;
assign enable_variable_to_check_86[2] = enable_variable_128_to_check_86;

// 拆分后校验节点86传递给变量节点166的值以及对变量节点166传递过来的值
wire [5:0] value_check_86_to_variable_166;
wire enable_check_86_to_variable_166;
wire [5:0] value_variable_166_to_check_86;
wire enable_variable_166_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_166 = value_check_86_to_variable[23:18];
assign enable_check_86_to_variable_166 = enable_check_86_to_variable[3];
// 对变量节点166传递过来的值进行组合
assign value_variable_to_check_86[23:18] = value_variable_166_to_check_86;
assign enable_variable_to_check_86[3] = enable_variable_166_to_check_86;

// 拆分后校验节点86传递给变量节点210的值以及对变量节点210传递过来的值
wire [5:0] value_check_86_to_variable_210;
wire enable_check_86_to_variable_210;
wire [5:0] value_variable_210_to_check_86;
wire enable_variable_210_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_210 = value_check_86_to_variable[29:24];
assign enable_check_86_to_variable_210 = enable_check_86_to_variable[4];
// 对变量节点210传递过来的值进行组合
assign value_variable_to_check_86[29:24] = value_variable_210_to_check_86;
assign enable_variable_to_check_86[4] = enable_variable_210_to_check_86;

// 拆分后校验节点86传递给变量节点232的值以及对变量节点232传递过来的值
wire [5:0] value_check_86_to_variable_232;
wire enable_check_86_to_variable_232;
wire [5:0] value_variable_232_to_check_86;
wire enable_variable_232_to_check_86;
// 对校验节点86的输出值进行拆分
assign value_check_86_to_variable_232 = value_check_86_to_variable[35:30];
assign enable_check_86_to_variable_232 = enable_check_86_to_variable[5];
// 对变量节点232传递过来的值进行组合
assign value_variable_to_check_86[35:30] = value_variable_232_to_check_86;
assign enable_variable_to_check_86[5] = enable_variable_232_to_check_86;


// 校验节点87的接口
wire [35:0] value_variable_to_check_87;
wire [35:0] value_check_87_to_variable;
wire [5:0] enable_variable_to_check_87;
wire [5:0] enable_check_87_to_variable;

// 拆分后校验节点87传递给变量节点29的值以及对变量节点29传递过来的值
wire [5:0] value_check_87_to_variable_29;
wire enable_check_87_to_variable_29;
wire [5:0] value_variable_29_to_check_87;
wire enable_variable_29_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_29 = value_check_87_to_variable[5:0];
assign enable_check_87_to_variable_29 = enable_check_87_to_variable[0];
// 对变量节点29传递过来的值进行组合
assign value_variable_to_check_87[5:0] = value_variable_29_to_check_87;
assign enable_variable_to_check_87[0] = enable_variable_29_to_check_87;

// 拆分后校验节点87传递给变量节点71的值以及对变量节点71传递过来的值
wire [5:0] value_check_87_to_variable_71;
wire enable_check_87_to_variable_71;
wire [5:0] value_variable_71_to_check_87;
wire enable_variable_71_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_71 = value_check_87_to_variable[11:6];
assign enable_check_87_to_variable_71 = enable_check_87_to_variable[1];
// 对变量节点71传递过来的值进行组合
assign value_variable_to_check_87[11:6] = value_variable_71_to_check_87;
assign enable_variable_to_check_87[1] = enable_variable_71_to_check_87;

// 拆分后校验节点87传递给变量节点98的值以及对变量节点98传递过来的值
wire [5:0] value_check_87_to_variable_98;
wire enable_check_87_to_variable_98;
wire [5:0] value_variable_98_to_check_87;
wire enable_variable_98_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_98 = value_check_87_to_variable[17:12];
assign enable_check_87_to_variable_98 = enable_check_87_to_variable[2];
// 对变量节点98传递过来的值进行组合
assign value_variable_to_check_87[17:12] = value_variable_98_to_check_87;
assign enable_variable_to_check_87[2] = enable_variable_98_to_check_87;

// 拆分后校验节点87传递给变量节点162的值以及对变量节点162传递过来的值
wire [5:0] value_check_87_to_variable_162;
wire enable_check_87_to_variable_162;
wire [5:0] value_variable_162_to_check_87;
wire enable_variable_162_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_162 = value_check_87_to_variable[23:18];
assign enable_check_87_to_variable_162 = enable_check_87_to_variable[3];
// 对变量节点162传递过来的值进行组合
assign value_variable_to_check_87[23:18] = value_variable_162_to_check_87;
assign enable_variable_to_check_87[3] = enable_variable_162_to_check_87;

// 拆分后校验节点87传递给变量节点208的值以及对变量节点208传递过来的值
wire [5:0] value_check_87_to_variable_208;
wire enable_check_87_to_variable_208;
wire [5:0] value_variable_208_to_check_87;
wire enable_variable_208_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_208 = value_check_87_to_variable[29:24];
assign enable_check_87_to_variable_208 = enable_check_87_to_variable[4];
// 对变量节点208传递过来的值进行组合
assign value_variable_to_check_87[29:24] = value_variable_208_to_check_87;
assign enable_variable_to_check_87[4] = enable_variable_208_to_check_87;

// 拆分后校验节点87传递给变量节点239的值以及对变量节点239传递过来的值
wire [5:0] value_check_87_to_variable_239;
wire enable_check_87_to_variable_239;
wire [5:0] value_variable_239_to_check_87;
wire enable_variable_239_to_check_87;
// 对校验节点87的输出值进行拆分
assign value_check_87_to_variable_239 = value_check_87_to_variable[35:30];
assign enable_check_87_to_variable_239 = enable_check_87_to_variable[5];
// 对变量节点239传递过来的值进行组合
assign value_variable_to_check_87[35:30] = value_variable_239_to_check_87;
assign enable_variable_to_check_87[5] = enable_variable_239_to_check_87;


// 校验节点88的接口
wire [35:0] value_variable_to_check_88;
wire [35:0] value_check_88_to_variable;
wire [5:0] enable_variable_to_check_88;
wire [5:0] enable_check_88_to_variable;

// 拆分后校验节点88传递给变量节点3的值以及对变量节点3传递过来的值
wire [5:0] value_check_88_to_variable_3;
wire enable_check_88_to_variable_3;
wire [5:0] value_variable_3_to_check_88;
wire enable_variable_3_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_3 = value_check_88_to_variable[5:0];
assign enable_check_88_to_variable_3 = enable_check_88_to_variable[0];
// 对变量节点3传递过来的值进行组合
assign value_variable_to_check_88[5:0] = value_variable_3_to_check_88;
assign enable_variable_to_check_88[0] = enable_variable_3_to_check_88;

// 拆分后校验节点88传递给变量节点52的值以及对变量节点52传递过来的值
wire [5:0] value_check_88_to_variable_52;
wire enable_check_88_to_variable_52;
wire [5:0] value_variable_52_to_check_88;
wire enable_variable_52_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_52 = value_check_88_to_variable[11:6];
assign enable_check_88_to_variable_52 = enable_check_88_to_variable[1];
// 对变量节点52传递过来的值进行组合
assign value_variable_to_check_88[11:6] = value_variable_52_to_check_88;
assign enable_variable_to_check_88[1] = enable_variable_52_to_check_88;

// 拆分后校验节点88传递给变量节点129的值以及对变量节点129传递过来的值
wire [5:0] value_check_88_to_variable_129;
wire enable_check_88_to_variable_129;
wire [5:0] value_variable_129_to_check_88;
wire enable_variable_129_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_129 = value_check_88_to_variable[17:12];
assign enable_check_88_to_variable_129 = enable_check_88_to_variable[2];
// 对变量节点129传递过来的值进行组合
assign value_variable_to_check_88[17:12] = value_variable_129_to_check_88;
assign enable_variable_to_check_88[2] = enable_variable_129_to_check_88;

// 拆分后校验节点88传递给变量节点167的值以及对变量节点167传递过来的值
wire [5:0] value_check_88_to_variable_167;
wire enable_check_88_to_variable_167;
wire [5:0] value_variable_167_to_check_88;
wire enable_variable_167_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_167 = value_check_88_to_variable[23:18];
assign enable_check_88_to_variable_167 = enable_check_88_to_variable[3];
// 对变量节点167传递过来的值进行组合
assign value_variable_to_check_88[23:18] = value_variable_167_to_check_88;
assign enable_variable_to_check_88[3] = enable_variable_167_to_check_88;

// 拆分后校验节点88传递给变量节点174的值以及对变量节点174传递过来的值
wire [5:0] value_check_88_to_variable_174;
wire enable_check_88_to_variable_174;
wire [5:0] value_variable_174_to_check_88;
wire enable_variable_174_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_174 = value_check_88_to_variable[29:24];
assign enable_check_88_to_variable_174 = enable_check_88_to_variable[4];
// 对变量节点174传递过来的值进行组合
assign value_variable_to_check_88[29:24] = value_variable_174_to_check_88;
assign enable_variable_to_check_88[4] = enable_variable_174_to_check_88;

// 拆分后校验节点88传递给变量节点247的值以及对变量节点247传递过来的值
wire [5:0] value_check_88_to_variable_247;
wire enable_check_88_to_variable_247;
wire [5:0] value_variable_247_to_check_88;
wire enable_variable_247_to_check_88;
// 对校验节点88的输出值进行拆分
assign value_check_88_to_variable_247 = value_check_88_to_variable[35:30];
assign enable_check_88_to_variable_247 = enable_check_88_to_variable[5];
// 对变量节点247传递过来的值进行组合
assign value_variable_to_check_88[35:30] = value_variable_247_to_check_88;
assign enable_variable_to_check_88[5] = enable_variable_247_to_check_88;


// 校验节点89的接口
wire [35:0] value_variable_to_check_89;
wire [35:0] value_check_89_to_variable;
wire [5:0] enable_variable_to_check_89;
wire [5:0] enable_check_89_to_variable;

// 拆分后校验节点89传递给变量节点37的值以及对变量节点37传递过来的值
wire [5:0] value_check_89_to_variable_37;
wire enable_check_89_to_variable_37;
wire [5:0] value_variable_37_to_check_89;
wire enable_variable_37_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_37 = value_check_89_to_variable[5:0];
assign enable_check_89_to_variable_37 = enable_check_89_to_variable[0];
// 对变量节点37传递过来的值进行组合
assign value_variable_to_check_89[5:0] = value_variable_37_to_check_89;
assign enable_variable_to_check_89[0] = enable_variable_37_to_check_89;

// 拆分后校验节点89传递给变量节点65的值以及对变量节点65传递过来的值
wire [5:0] value_check_89_to_variable_65;
wire enable_check_89_to_variable_65;
wire [5:0] value_variable_65_to_check_89;
wire enable_variable_65_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_65 = value_check_89_to_variable[11:6];
assign enable_check_89_to_variable_65 = enable_check_89_to_variable[1];
// 对变量节点65传递过来的值进行组合
assign value_variable_to_check_89[11:6] = value_variable_65_to_check_89;
assign enable_variable_to_check_89[1] = enable_variable_65_to_check_89;

// 拆分后校验节点89传递给变量节点122的值以及对变量节点122传递过来的值
wire [5:0] value_check_89_to_variable_122;
wire enable_check_89_to_variable_122;
wire [5:0] value_variable_122_to_check_89;
wire enable_variable_122_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_122 = value_check_89_to_variable[17:12];
assign enable_check_89_to_variable_122 = enable_check_89_to_variable[2];
// 对变量节点122传递过来的值进行组合
assign value_variable_to_check_89[17:12] = value_variable_122_to_check_89;
assign enable_variable_to_check_89[2] = enable_variable_122_to_check_89;

// 拆分后校验节点89传递给变量节点147的值以及对变量节点147传递过来的值
wire [5:0] value_check_89_to_variable_147;
wire enable_check_89_to_variable_147;
wire [5:0] value_variable_147_to_check_89;
wire enable_variable_147_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_147 = value_check_89_to_variable[23:18];
assign enable_check_89_to_variable_147 = enable_check_89_to_variable[3];
// 对变量节点147传递过来的值进行组合
assign value_variable_to_check_89[23:18] = value_variable_147_to_check_89;
assign enable_variable_to_check_89[3] = enable_variable_147_to_check_89;

// 拆分后校验节点89传递给变量节点196的值以及对变量节点196传递过来的值
wire [5:0] value_check_89_to_variable_196;
wire enable_check_89_to_variable_196;
wire [5:0] value_variable_196_to_check_89;
wire enable_variable_196_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_196 = value_check_89_to_variable[29:24];
assign enable_check_89_to_variable_196 = enable_check_89_to_variable[4];
// 对变量节点196传递过来的值进行组合
assign value_variable_to_check_89[29:24] = value_variable_196_to_check_89;
assign enable_variable_to_check_89[4] = enable_variable_196_to_check_89;

// 拆分后校验节点89传递给变量节点219的值以及对变量节点219传递过来的值
wire [5:0] value_check_89_to_variable_219;
wire enable_check_89_to_variable_219;
wire [5:0] value_variable_219_to_check_89;
wire enable_variable_219_to_check_89;
// 对校验节点89的输出值进行拆分
assign value_check_89_to_variable_219 = value_check_89_to_variable[35:30];
assign enable_check_89_to_variable_219 = enable_check_89_to_variable[5];
// 对变量节点219传递过来的值进行组合
assign value_variable_to_check_89[35:30] = value_variable_219_to_check_89;
assign enable_variable_to_check_89[5] = enable_variable_219_to_check_89;


// 校验节点90的接口
wire [35:0] value_variable_to_check_90;
wire [35:0] value_check_90_to_variable;
wire [5:0] enable_variable_to_check_90;
wire [5:0] enable_check_90_to_variable;

// 拆分后校验节点90传递给变量节点14的值以及对变量节点14传递过来的值
wire [5:0] value_check_90_to_variable_14;
wire enable_check_90_to_variable_14;
wire [5:0] value_variable_14_to_check_90;
wire enable_variable_14_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_14 = value_check_90_to_variable[5:0];
assign enable_check_90_to_variable_14 = enable_check_90_to_variable[0];
// 对变量节点14传递过来的值进行组合
assign value_variable_to_check_90[5:0] = value_variable_14_to_check_90;
assign enable_variable_to_check_90[0] = enable_variable_14_to_check_90;

// 拆分后校验节点90传递给变量节点82的值以及对变量节点82传递过来的值
wire [5:0] value_check_90_to_variable_82;
wire enable_check_90_to_variable_82;
wire [5:0] value_variable_82_to_check_90;
wire enable_variable_82_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_82 = value_check_90_to_variable[11:6];
assign enable_check_90_to_variable_82 = enable_check_90_to_variable[1];
// 对变量节点82传递过来的值进行组合
assign value_variable_to_check_90[11:6] = value_variable_82_to_check_90;
assign enable_variable_to_check_90[1] = enable_variable_82_to_check_90;

// 拆分后校验节点90传递给变量节点112的值以及对变量节点112传递过来的值
wire [5:0] value_check_90_to_variable_112;
wire enable_check_90_to_variable_112;
wire [5:0] value_variable_112_to_check_90;
wire enable_variable_112_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_112 = value_check_90_to_variable[17:12];
assign enable_check_90_to_variable_112 = enable_check_90_to_variable[2];
// 对变量节点112传递过来的值进行组合
assign value_variable_to_check_90[17:12] = value_variable_112_to_check_90;
assign enable_variable_to_check_90[2] = enable_variable_112_to_check_90;

// 拆分后校验节点90传递给变量节点137的值以及对变量节点137传递过来的值
wire [5:0] value_check_90_to_variable_137;
wire enable_check_90_to_variable_137;
wire [5:0] value_variable_137_to_check_90;
wire enable_variable_137_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_137 = value_check_90_to_variable[23:18];
assign enable_check_90_to_variable_137 = enable_check_90_to_variable[3];
// 对变量节点137传递过来的值进行组合
assign value_variable_to_check_90[23:18] = value_variable_137_to_check_90;
assign enable_variable_to_check_90[3] = enable_variable_137_to_check_90;

// 拆分后校验节点90传递给变量节点207的值以及对变量节点207传递过来的值
wire [5:0] value_check_90_to_variable_207;
wire enable_check_90_to_variable_207;
wire [5:0] value_variable_207_to_check_90;
wire enable_variable_207_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_207 = value_check_90_to_variable[29:24];
assign enable_check_90_to_variable_207 = enable_check_90_to_variable[4];
// 对变量节点207传递过来的值进行组合
assign value_variable_to_check_90[29:24] = value_variable_207_to_check_90;
assign enable_variable_to_check_90[4] = enable_variable_207_to_check_90;

// 拆分后校验节点90传递给变量节点246的值以及对变量节点246传递过来的值
wire [5:0] value_check_90_to_variable_246;
wire enable_check_90_to_variable_246;
wire [5:0] value_variable_246_to_check_90;
wire enable_variable_246_to_check_90;
// 对校验节点90的输出值进行拆分
assign value_check_90_to_variable_246 = value_check_90_to_variable[35:30];
assign enable_check_90_to_variable_246 = enable_check_90_to_variable[5];
// 对变量节点246传递过来的值进行组合
assign value_variable_to_check_90[35:30] = value_variable_246_to_check_90;
assign enable_variable_to_check_90[5] = enable_variable_246_to_check_90;


// 校验节点91的接口
wire [35:0] value_variable_to_check_91;
wire [35:0] value_check_91_to_variable;
wire [5:0] enable_variable_to_check_91;
wire [5:0] enable_check_91_to_variable;

// 拆分后校验节点91传递给变量节点4的值以及对变量节点4传递过来的值
wire [5:0] value_check_91_to_variable_4;
wire enable_check_91_to_variable_4;
wire [5:0] value_variable_4_to_check_91;
wire enable_variable_4_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_4 = value_check_91_to_variable[5:0];
assign enable_check_91_to_variable_4 = enable_check_91_to_variable[0];
// 对变量节点4传递过来的值进行组合
assign value_variable_to_check_91[5:0] = value_variable_4_to_check_91;
assign enable_variable_to_check_91[0] = enable_variable_4_to_check_91;

// 拆分后校验节点91传递给变量节点71的值以及对变量节点71传递过来的值
wire [5:0] value_check_91_to_variable_71;
wire enable_check_91_to_variable_71;
wire [5:0] value_variable_71_to_check_91;
wire enable_variable_71_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_71 = value_check_91_to_variable[11:6];
assign enable_check_91_to_variable_71 = enable_check_91_to_variable[1];
// 对变量节点71传递过来的值进行组合
assign value_variable_to_check_91[11:6] = value_variable_71_to_check_91;
assign enable_variable_to_check_91[1] = enable_variable_71_to_check_91;

// 拆分后校验节点91传递给变量节点121的值以及对变量节点121传递过来的值
wire [5:0] value_check_91_to_variable_121;
wire enable_check_91_to_variable_121;
wire [5:0] value_variable_121_to_check_91;
wire enable_variable_121_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_121 = value_check_91_to_variable[17:12];
assign enable_check_91_to_variable_121 = enable_check_91_to_variable[2];
// 对变量节点121传递过来的值进行组合
assign value_variable_to_check_91[17:12] = value_variable_121_to_check_91;
assign enable_variable_to_check_91[2] = enable_variable_121_to_check_91;

// 拆分后校验节点91传递给变量节点161的值以及对变量节点161传递过来的值
wire [5:0] value_check_91_to_variable_161;
wire enable_check_91_to_variable_161;
wire [5:0] value_variable_161_to_check_91;
wire enable_variable_161_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_161 = value_check_91_to_variable[23:18];
assign enable_check_91_to_variable_161 = enable_check_91_to_variable[3];
// 对变量节点161传递过来的值进行组合
assign value_variable_to_check_91[23:18] = value_variable_161_to_check_91;
assign enable_variable_to_check_91[3] = enable_variable_161_to_check_91;

// 拆分后校验节点91传递给变量节点190的值以及对变量节点190传递过来的值
wire [5:0] value_check_91_to_variable_190;
wire enable_check_91_to_variable_190;
wire [5:0] value_variable_190_to_check_91;
wire enable_variable_190_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_190 = value_check_91_to_variable[29:24];
assign enable_check_91_to_variable_190 = enable_check_91_to_variable[4];
// 对变量节点190传递过来的值进行组合
assign value_variable_to_check_91[29:24] = value_variable_190_to_check_91;
assign enable_variable_to_check_91[4] = enable_variable_190_to_check_91;

// 拆分后校验节点91传递给变量节点230的值以及对变量节点230传递过来的值
wire [5:0] value_check_91_to_variable_230;
wire enable_check_91_to_variable_230;
wire [5:0] value_variable_230_to_check_91;
wire enable_variable_230_to_check_91;
// 对校验节点91的输出值进行拆分
assign value_check_91_to_variable_230 = value_check_91_to_variable[35:30];
assign enable_check_91_to_variable_230 = enable_check_91_to_variable[5];
// 对变量节点230传递过来的值进行组合
assign value_variable_to_check_91[35:30] = value_variable_230_to_check_91;
assign enable_variable_to_check_91[5] = enable_variable_230_to_check_91;


// 校验节点92的接口
wire [35:0] value_variable_to_check_92;
wire [35:0] value_check_92_to_variable;
wire [5:0] enable_variable_to_check_92;
wire [5:0] enable_check_92_to_variable;

// 拆分后校验节点92传递给变量节点40的值以及对变量节点40传递过来的值
wire [5:0] value_check_92_to_variable_40;
wire enable_check_92_to_variable_40;
wire [5:0] value_variable_40_to_check_92;
wire enable_variable_40_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_40 = value_check_92_to_variable[5:0];
assign enable_check_92_to_variable_40 = enable_check_92_to_variable[0];
// 对变量节点40传递过来的值进行组合
assign value_variable_to_check_92[5:0] = value_variable_40_to_check_92;
assign enable_variable_to_check_92[0] = enable_variable_40_to_check_92;

// 拆分后校验节点92传递给变量节点70的值以及对变量节点70传递过来的值
wire [5:0] value_check_92_to_variable_70;
wire enable_check_92_to_variable_70;
wire [5:0] value_variable_70_to_check_92;
wire enable_variable_70_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_70 = value_check_92_to_variable[11:6];
assign enable_check_92_to_variable_70 = enable_check_92_to_variable[1];
// 对变量节点70传递过来的值进行组合
assign value_variable_to_check_92[11:6] = value_variable_70_to_check_92;
assign enable_variable_to_check_92[1] = enable_variable_70_to_check_92;

// 拆分后校验节点92传递给变量节点108的值以及对变量节点108传递过来的值
wire [5:0] value_check_92_to_variable_108;
wire enable_check_92_to_variable_108;
wire [5:0] value_variable_108_to_check_92;
wire enable_variable_108_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_108 = value_check_92_to_variable[17:12];
assign enable_check_92_to_variable_108 = enable_check_92_to_variable[2];
// 对变量节点108传递过来的值进行组合
assign value_variable_to_check_92[17:12] = value_variable_108_to_check_92;
assign enable_variable_to_check_92[2] = enable_variable_108_to_check_92;

// 拆分后校验节点92传递给变量节点133的值以及对变量节点133传递过来的值
wire [5:0] value_check_92_to_variable_133;
wire enable_check_92_to_variable_133;
wire [5:0] value_variable_133_to_check_92;
wire enable_variable_133_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_133 = value_check_92_to_variable[23:18];
assign enable_check_92_to_variable_133 = enable_check_92_to_variable[3];
// 对变量节点133传递过来的值进行组合
assign value_variable_to_check_92[23:18] = value_variable_133_to_check_92;
assign enable_variable_to_check_92[3] = enable_variable_133_to_check_92;

// 拆分后校验节点92传递给变量节点207的值以及对变量节点207传递过来的值
wire [5:0] value_check_92_to_variable_207;
wire enable_check_92_to_variable_207;
wire [5:0] value_variable_207_to_check_92;
wire enable_variable_207_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_207 = value_check_92_to_variable[29:24];
assign enable_check_92_to_variable_207 = enable_check_92_to_variable[4];
// 对变量节点207传递过来的值进行组合
assign value_variable_to_check_92[29:24] = value_variable_207_to_check_92;
assign enable_variable_to_check_92[4] = enable_variable_207_to_check_92;

// 拆分后校验节点92传递给变量节点226的值以及对变量节点226传递过来的值
wire [5:0] value_check_92_to_variable_226;
wire enable_check_92_to_variable_226;
wire [5:0] value_variable_226_to_check_92;
wire enable_variable_226_to_check_92;
// 对校验节点92的输出值进行拆分
assign value_check_92_to_variable_226 = value_check_92_to_variable[35:30];
assign enable_check_92_to_variable_226 = enable_check_92_to_variable[5];
// 对变量节点226传递过来的值进行组合
assign value_variable_to_check_92[35:30] = value_variable_226_to_check_92;
assign enable_variable_to_check_92[5] = enable_variable_226_to_check_92;


// 校验节点93的接口
wire [35:0] value_variable_to_check_93;
wire [35:0] value_check_93_to_variable;
wire [5:0] enable_variable_to_check_93;
wire [5:0] enable_check_93_to_variable;

// 拆分后校验节点93传递给变量节点8的值以及对变量节点8传递过来的值
wire [5:0] value_check_93_to_variable_8;
wire enable_check_93_to_variable_8;
wire [5:0] value_variable_8_to_check_93;
wire enable_variable_8_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_8 = value_check_93_to_variable[5:0];
assign enable_check_93_to_variable_8 = enable_check_93_to_variable[0];
// 对变量节点8传递过来的值进行组合
assign value_variable_to_check_93[5:0] = value_variable_8_to_check_93;
assign enable_variable_to_check_93[0] = enable_variable_8_to_check_93;

// 拆分后校验节点93传递给变量节点72的值以及对变量节点72传递过来的值
wire [5:0] value_check_93_to_variable_72;
wire enable_check_93_to_variable_72;
wire [5:0] value_variable_72_to_check_93;
wire enable_variable_72_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_72 = value_check_93_to_variable[11:6];
assign enable_check_93_to_variable_72 = enable_check_93_to_variable[1];
// 对变量节点72传递过来的值进行组合
assign value_variable_to_check_93[11:6] = value_variable_72_to_check_93;
assign enable_variable_to_check_93[1] = enable_variable_72_to_check_93;

// 拆分后校验节点93传递给变量节点118的值以及对变量节点118传递过来的值
wire [5:0] value_check_93_to_variable_118;
wire enable_check_93_to_variable_118;
wire [5:0] value_variable_118_to_check_93;
wire enable_variable_118_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_118 = value_check_93_to_variable[17:12];
assign enable_check_93_to_variable_118 = enable_check_93_to_variable[2];
// 对变量节点118传递过来的值进行组合
assign value_variable_to_check_93[17:12] = value_variable_118_to_check_93;
assign enable_variable_to_check_93[2] = enable_variable_118_to_check_93;

// 拆分后校验节点93传递给变量节点161的值以及对变量节点161传递过来的值
wire [5:0] value_check_93_to_variable_161;
wire enable_check_93_to_variable_161;
wire [5:0] value_variable_161_to_check_93;
wire enable_variable_161_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_161 = value_check_93_to_variable[23:18];
assign enable_check_93_to_variable_161 = enable_check_93_to_variable[3];
// 对变量节点161传递过来的值进行组合
assign value_variable_to_check_93[23:18] = value_variable_161_to_check_93;
assign enable_variable_to_check_93[3] = enable_variable_161_to_check_93;

// 拆分后校验节点93传递给变量节点199的值以及对变量节点199传递过来的值
wire [5:0] value_check_93_to_variable_199;
wire enable_check_93_to_variable_199;
wire [5:0] value_variable_199_to_check_93;
wire enable_variable_199_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_199 = value_check_93_to_variable[29:24];
assign enable_check_93_to_variable_199 = enable_check_93_to_variable[4];
// 对变量节点199传递过来的值进行组合
assign value_variable_to_check_93[29:24] = value_variable_199_to_check_93;
assign enable_variable_to_check_93[4] = enable_variable_199_to_check_93;

// 拆分后校验节点93传递给变量节点247的值以及对变量节点247传递过来的值
wire [5:0] value_check_93_to_variable_247;
wire enable_check_93_to_variable_247;
wire [5:0] value_variable_247_to_check_93;
wire enable_variable_247_to_check_93;
// 对校验节点93的输出值进行拆分
assign value_check_93_to_variable_247 = value_check_93_to_variable[35:30];
assign enable_check_93_to_variable_247 = enable_check_93_to_variable[5];
// 对变量节点247传递过来的值进行组合
assign value_variable_to_check_93[35:30] = value_variable_247_to_check_93;
assign enable_variable_to_check_93[5] = enable_variable_247_to_check_93;


// 校验节点94的接口
wire [35:0] value_variable_to_check_94;
wire [35:0] value_check_94_to_variable;
wire [5:0] enable_variable_to_check_94;
wire [5:0] enable_check_94_to_variable;

// 拆分后校验节点94传递给变量节点9的值以及对变量节点9传递过来的值
wire [5:0] value_check_94_to_variable_9;
wire enable_check_94_to_variable_9;
wire [5:0] value_variable_9_to_check_94;
wire enable_variable_9_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_9 = value_check_94_to_variable[5:0];
assign enable_check_94_to_variable_9 = enable_check_94_to_variable[0];
// 对变量节点9传递过来的值进行组合
assign value_variable_to_check_94[5:0] = value_variable_9_to_check_94;
assign enable_variable_to_check_94[0] = enable_variable_9_to_check_94;

// 拆分后校验节点94传递给变量节点79的值以及对变量节点79传递过来的值
wire [5:0] value_check_94_to_variable_79;
wire enable_check_94_to_variable_79;
wire [5:0] value_variable_79_to_check_94;
wire enable_variable_79_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_79 = value_check_94_to_variable[11:6];
assign enable_check_94_to_variable_79 = enable_check_94_to_variable[1];
// 对变量节点79传递过来的值进行组合
assign value_variable_to_check_94[11:6] = value_variable_79_to_check_94;
assign enable_variable_to_check_94[1] = enable_variable_79_to_check_94;

// 拆分后校验节点94传递给变量节点120的值以及对变量节点120传递过来的值
wire [5:0] value_check_94_to_variable_120;
wire enable_check_94_to_variable_120;
wire [5:0] value_variable_120_to_check_94;
wire enable_variable_120_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_120 = value_check_94_to_variable[17:12];
assign enable_check_94_to_variable_120 = enable_check_94_to_variable[2];
// 对变量节点120传递过来的值进行组合
assign value_variable_to_check_94[17:12] = value_variable_120_to_check_94;
assign enable_variable_to_check_94[2] = enable_variable_120_to_check_94;

// 拆分后校验节点94传递给变量节点133的值以及对变量节点133传递过来的值
wire [5:0] value_check_94_to_variable_133;
wire enable_check_94_to_variable_133;
wire [5:0] value_variable_133_to_check_94;
wire enable_variable_133_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_133 = value_check_94_to_variable[23:18];
assign enable_check_94_to_variable_133 = enable_check_94_to_variable[3];
// 对变量节点133传递过来的值进行组合
assign value_variable_to_check_94[23:18] = value_variable_133_to_check_94;
assign enable_variable_to_check_94[3] = enable_variable_133_to_check_94;

// 拆分后校验节点94传递给变量节点192的值以及对变量节点192传递过来的值
wire [5:0] value_check_94_to_variable_192;
wire enable_check_94_to_variable_192;
wire [5:0] value_variable_192_to_check_94;
wire enable_variable_192_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_192 = value_check_94_to_variable[29:24];
assign enable_check_94_to_variable_192 = enable_check_94_to_variable[4];
// 对变量节点192传递过来的值进行组合
assign value_variable_to_check_94[29:24] = value_variable_192_to_check_94;
assign enable_variable_to_check_94[4] = enable_variable_192_to_check_94;

// 拆分后校验节点94传递给变量节点244的值以及对变量节点244传递过来的值
wire [5:0] value_check_94_to_variable_244;
wire enable_check_94_to_variable_244;
wire [5:0] value_variable_244_to_check_94;
wire enable_variable_244_to_check_94;
// 对校验节点94的输出值进行拆分
assign value_check_94_to_variable_244 = value_check_94_to_variable[35:30];
assign enable_check_94_to_variable_244 = enable_check_94_to_variable[5];
// 对变量节点244传递过来的值进行组合
assign value_variable_to_check_94[35:30] = value_variable_244_to_check_94;
assign enable_variable_to_check_94[5] = enable_variable_244_to_check_94;


// 校验节点95的接口
wire [35:0] value_variable_to_check_95;
wire [35:0] value_check_95_to_variable;
wire [5:0] enable_variable_to_check_95;
wire [5:0] enable_check_95_to_variable;

// 拆分后校验节点95传递给变量节点16的值以及对变量节点16传递过来的值
wire [5:0] value_check_95_to_variable_16;
wire enable_check_95_to_variable_16;
wire [5:0] value_variable_16_to_check_95;
wire enable_variable_16_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_16 = value_check_95_to_variable[5:0];
assign enable_check_95_to_variable_16 = enable_check_95_to_variable[0];
// 对变量节点16传递过来的值进行组合
assign value_variable_to_check_95[5:0] = value_variable_16_to_check_95;
assign enable_variable_to_check_95[0] = enable_variable_16_to_check_95;

// 拆分后校验节点95传递给变量节点59的值以及对变量节点59传递过来的值
wire [5:0] value_check_95_to_variable_59;
wire enable_check_95_to_variable_59;
wire [5:0] value_variable_59_to_check_95;
wire enable_variable_59_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_59 = value_check_95_to_variable[11:6];
assign enable_check_95_to_variable_59 = enable_check_95_to_variable[1];
// 对变量节点59传递过来的值进行组合
assign value_variable_to_check_95[11:6] = value_variable_59_to_check_95;
assign enable_variable_to_check_95[1] = enable_variable_59_to_check_95;

// 拆分后校验节点95传递给变量节点124的值以及对变量节点124传递过来的值
wire [5:0] value_check_95_to_variable_124;
wire enable_check_95_to_variable_124;
wire [5:0] value_variable_124_to_check_95;
wire enable_variable_124_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_124 = value_check_95_to_variable[17:12];
assign enable_check_95_to_variable_124 = enable_check_95_to_variable[2];
// 对变量节点124传递过来的值进行组合
assign value_variable_to_check_95[17:12] = value_variable_124_to_check_95;
assign enable_variable_to_check_95[2] = enable_variable_124_to_check_95;

// 拆分后校验节点95传递给变量节点168的值以及对变量节点168传递过来的值
wire [5:0] value_check_95_to_variable_168;
wire enable_check_95_to_variable_168;
wire [5:0] value_variable_168_to_check_95;
wire enable_variable_168_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_168 = value_check_95_to_variable[23:18];
assign enable_check_95_to_variable_168 = enable_check_95_to_variable[3];
// 对变量节点168传递过来的值进行组合
assign value_variable_to_check_95[23:18] = value_variable_168_to_check_95;
assign enable_variable_to_check_95[3] = enable_variable_168_to_check_95;

// 拆分后校验节点95传递给变量节点208的值以及对变量节点208传递过来的值
wire [5:0] value_check_95_to_variable_208;
wire enable_check_95_to_variable_208;
wire [5:0] value_variable_208_to_check_95;
wire enable_variable_208_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_208 = value_check_95_to_variable[29:24];
assign enable_check_95_to_variable_208 = enable_check_95_to_variable[4];
// 对变量节点208传递过来的值进行组合
assign value_variable_to_check_95[29:24] = value_variable_208_to_check_95;
assign enable_variable_to_check_95[4] = enable_variable_208_to_check_95;

// 拆分后校验节点95传递给变量节点255的值以及对变量节点255传递过来的值
wire [5:0] value_check_95_to_variable_255;
wire enable_check_95_to_variable_255;
wire [5:0] value_variable_255_to_check_95;
wire enable_variable_255_to_check_95;
// 对校验节点95的输出值进行拆分
assign value_check_95_to_variable_255 = value_check_95_to_variable[35:30];
assign enable_check_95_to_variable_255 = enable_check_95_to_variable[5];
// 对变量节点255传递过来的值进行组合
assign value_variable_to_check_95[35:30] = value_variable_255_to_check_95;
assign enable_variable_to_check_95[5] = enable_variable_255_to_check_95;


// 校验节点96的接口
wire [35:0] value_variable_to_check_96;
wire [35:0] value_check_96_to_variable;
wire [5:0] enable_variable_to_check_96;
wire [5:0] enable_check_96_to_variable;

// 拆分后校验节点96传递给变量节点13的值以及对变量节点13传递过来的值
wire [5:0] value_check_96_to_variable_13;
wire enable_check_96_to_variable_13;
wire [5:0] value_variable_13_to_check_96;
wire enable_variable_13_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_13 = value_check_96_to_variable[5:0];
assign enable_check_96_to_variable_13 = enable_check_96_to_variable[0];
// 对变量节点13传递过来的值进行组合
assign value_variable_to_check_96[5:0] = value_variable_13_to_check_96;
assign enable_variable_to_check_96[0] = enable_variable_13_to_check_96;

// 拆分后校验节点96传递给变量节点45的值以及对变量节点45传递过来的值
wire [5:0] value_check_96_to_variable_45;
wire enable_check_96_to_variable_45;
wire [5:0] value_variable_45_to_check_96;
wire enable_variable_45_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_45 = value_check_96_to_variable[11:6];
assign enable_check_96_to_variable_45 = enable_check_96_to_variable[1];
// 对变量节点45传递过来的值进行组合
assign value_variable_to_check_96[11:6] = value_variable_45_to_check_96;
assign enable_variable_to_check_96[1] = enable_variable_45_to_check_96;

// 拆分后校验节点96传递给变量节点128的值以及对变量节点128传递过来的值
wire [5:0] value_check_96_to_variable_128;
wire enable_check_96_to_variable_128;
wire [5:0] value_variable_128_to_check_96;
wire enable_variable_128_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_128 = value_check_96_to_variable[17:12];
assign enable_check_96_to_variable_128 = enable_check_96_to_variable[2];
// 对变量节点128传递过来的值进行组合
assign value_variable_to_check_96[17:12] = value_variable_128_to_check_96;
assign enable_variable_to_check_96[2] = enable_variable_128_to_check_96;

// 拆分后校验节点96传递给变量节点151的值以及对变量节点151传递过来的值
wire [5:0] value_check_96_to_variable_151;
wire enable_check_96_to_variable_151;
wire [5:0] value_variable_151_to_check_96;
wire enable_variable_151_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_151 = value_check_96_to_variable[23:18];
assign enable_check_96_to_variable_151 = enable_check_96_to_variable[3];
// 对变量节点151传递过来的值进行组合
assign value_variable_to_check_96[23:18] = value_variable_151_to_check_96;
assign enable_variable_to_check_96[3] = enable_variable_151_to_check_96;

// 拆分后校验节点96传递给变量节点178的值以及对变量节点178传递过来的值
wire [5:0] value_check_96_to_variable_178;
wire enable_check_96_to_variable_178;
wire [5:0] value_variable_178_to_check_96;
wire enable_variable_178_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_178 = value_check_96_to_variable[29:24];
assign enable_check_96_to_variable_178 = enable_check_96_to_variable[4];
// 对变量节点178传递过来的值进行组合
assign value_variable_to_check_96[29:24] = value_variable_178_to_check_96;
assign enable_variable_to_check_96[4] = enable_variable_178_to_check_96;

// 拆分后校验节点96传递给变量节点250的值以及对变量节点250传递过来的值
wire [5:0] value_check_96_to_variable_250;
wire enable_check_96_to_variable_250;
wire [5:0] value_variable_250_to_check_96;
wire enable_variable_250_to_check_96;
// 对校验节点96的输出值进行拆分
assign value_check_96_to_variable_250 = value_check_96_to_variable[35:30];
assign enable_check_96_to_variable_250 = enable_check_96_to_variable[5];
// 对变量节点250传递过来的值进行组合
assign value_variable_to_check_96[35:30] = value_variable_250_to_check_96;
assign enable_variable_to_check_96[5] = enable_variable_250_to_check_96;


// 校验节点97的接口
wire [35:0] value_variable_to_check_97;
wire [35:0] value_check_97_to_variable;
wire [5:0] enable_variable_to_check_97;
wire [5:0] enable_check_97_to_variable;

// 拆分后校验节点97传递给变量节点41的值以及对变量节点41传递过来的值
wire [5:0] value_check_97_to_variable_41;
wire enable_check_97_to_variable_41;
wire [5:0] value_variable_41_to_check_97;
wire enable_variable_41_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_41 = value_check_97_to_variable[5:0];
assign enable_check_97_to_variable_41 = enable_check_97_to_variable[0];
// 对变量节点41传递过来的值进行组合
assign value_variable_to_check_97[5:0] = value_variable_41_to_check_97;
assign enable_variable_to_check_97[0] = enable_variable_41_to_check_97;

// 拆分后校验节点97传递给变量节点54的值以及对变量节点54传递过来的值
wire [5:0] value_check_97_to_variable_54;
wire enable_check_97_to_variable_54;
wire [5:0] value_variable_54_to_check_97;
wire enable_variable_54_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_54 = value_check_97_to_variable[11:6];
assign enable_check_97_to_variable_54 = enable_check_97_to_variable[1];
// 对变量节点54传递过来的值进行组合
assign value_variable_to_check_97[11:6] = value_variable_54_to_check_97;
assign enable_variable_to_check_97[1] = enable_variable_54_to_check_97;

// 拆分后校验节点97传递给变量节点88的值以及对变量节点88传递过来的值
wire [5:0] value_check_97_to_variable_88;
wire enable_check_97_to_variable_88;
wire [5:0] value_variable_88_to_check_97;
wire enable_variable_88_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_88 = value_check_97_to_variable[17:12];
assign enable_check_97_to_variable_88 = enable_check_97_to_variable[2];
// 对变量节点88传递过来的值进行组合
assign value_variable_to_check_97[17:12] = value_variable_88_to_check_97;
assign enable_variable_to_check_97[2] = enable_variable_88_to_check_97;

// 拆分后校验节点97传递给变量节点149的值以及对变量节点149传递过来的值
wire [5:0] value_check_97_to_variable_149;
wire enable_check_97_to_variable_149;
wire [5:0] value_variable_149_to_check_97;
wire enable_variable_149_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_149 = value_check_97_to_variable[23:18];
assign enable_check_97_to_variable_149 = enable_check_97_to_variable[3];
// 对变量节点149传递过来的值进行组合
assign value_variable_to_check_97[23:18] = value_variable_149_to_check_97;
assign enable_variable_to_check_97[3] = enable_variable_149_to_check_97;

// 拆分后校验节点97传递给变量节点211的值以及对变量节点211传递过来的值
wire [5:0] value_check_97_to_variable_211;
wire enable_check_97_to_variable_211;
wire [5:0] value_variable_211_to_check_97;
wire enable_variable_211_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_211 = value_check_97_to_variable[29:24];
assign enable_check_97_to_variable_211 = enable_check_97_to_variable[4];
// 对变量节点211传递过来的值进行组合
assign value_variable_to_check_97[29:24] = value_variable_211_to_check_97;
assign enable_variable_to_check_97[4] = enable_variable_211_to_check_97;

// 拆分后校验节点97传递给变量节点240的值以及对变量节点240传递过来的值
wire [5:0] value_check_97_to_variable_240;
wire enable_check_97_to_variable_240;
wire [5:0] value_variable_240_to_check_97;
wire enable_variable_240_to_check_97;
// 对校验节点97的输出值进行拆分
assign value_check_97_to_variable_240 = value_check_97_to_variable[35:30];
assign enable_check_97_to_variable_240 = enable_check_97_to_variable[5];
// 对变量节点240传递过来的值进行组合
assign value_variable_to_check_97[35:30] = value_variable_240_to_check_97;
assign enable_variable_to_check_97[5] = enable_variable_240_to_check_97;


// 校验节点98的接口
wire [35:0] value_variable_to_check_98;
wire [35:0] value_check_98_to_variable;
wire [5:0] enable_variable_to_check_98;
wire [5:0] enable_check_98_to_variable;

// 拆分后校验节点98传递给变量节点34的值以及对变量节点34传递过来的值
wire [5:0] value_check_98_to_variable_34;
wire enable_check_98_to_variable_34;
wire [5:0] value_variable_34_to_check_98;
wire enable_variable_34_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_34 = value_check_98_to_variable[5:0];
assign enable_check_98_to_variable_34 = enable_check_98_to_variable[0];
// 对变量节点34传递过来的值进行组合
assign value_variable_to_check_98[5:0] = value_variable_34_to_check_98;
assign enable_variable_to_check_98[0] = enable_variable_34_to_check_98;

// 拆分后校验节点98传递给变量节点67的值以及对变量节点67传递过来的值
wire [5:0] value_check_98_to_variable_67;
wire enable_check_98_to_variable_67;
wire [5:0] value_variable_67_to_check_98;
wire enable_variable_67_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_67 = value_check_98_to_variable[11:6];
assign enable_check_98_to_variable_67 = enable_check_98_to_variable[1];
// 对变量节点67传递过来的值进行组合
assign value_variable_to_check_98[11:6] = value_variable_67_to_check_98;
assign enable_variable_to_check_98[1] = enable_variable_67_to_check_98;

// 拆分后校验节点98传递给变量节点95的值以及对变量节点95传递过来的值
wire [5:0] value_check_98_to_variable_95;
wire enable_check_98_to_variable_95;
wire [5:0] value_variable_95_to_check_98;
wire enable_variable_95_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_95 = value_check_98_to_variable[17:12];
assign enable_check_98_to_variable_95 = enable_check_98_to_variable[2];
// 对变量节点95传递过来的值进行组合
assign value_variable_to_check_98[17:12] = value_variable_95_to_check_98;
assign enable_variable_to_check_98[2] = enable_variable_95_to_check_98;

// 拆分后校验节点98传递给变量节点169的值以及对变量节点169传递过来的值
wire [5:0] value_check_98_to_variable_169;
wire enable_check_98_to_variable_169;
wire [5:0] value_variable_169_to_check_98;
wire enable_variable_169_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_169 = value_check_98_to_variable[23:18];
assign enable_check_98_to_variable_169 = enable_check_98_to_variable[3];
// 对变量节点169传递过来的值进行组合
assign value_variable_to_check_98[23:18] = value_variable_169_to_check_98;
assign enable_variable_to_check_98[3] = enable_variable_169_to_check_98;

// 拆分后校验节点98传递给变量节点173的值以及对变量节点173传递过来的值
wire [5:0] value_check_98_to_variable_173;
wire enable_check_98_to_variable_173;
wire [5:0] value_variable_173_to_check_98;
wire enable_variable_173_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_173 = value_check_98_to_variable[29:24];
assign enable_check_98_to_variable_173 = enable_check_98_to_variable[4];
// 对变量节点173传递过来的值进行组合
assign value_variable_to_check_98[29:24] = value_variable_173_to_check_98;
assign enable_variable_to_check_98[4] = enable_variable_173_to_check_98;

// 拆分后校验节点98传递给变量节点233的值以及对变量节点233传递过来的值
wire [5:0] value_check_98_to_variable_233;
wire enable_check_98_to_variable_233;
wire [5:0] value_variable_233_to_check_98;
wire enable_variable_233_to_check_98;
// 对校验节点98的输出值进行拆分
assign value_check_98_to_variable_233 = value_check_98_to_variable[35:30];
assign enable_check_98_to_variable_233 = enable_check_98_to_variable[5];
// 对变量节点233传递过来的值进行组合
assign value_variable_to_check_98[35:30] = value_variable_233_to_check_98;
assign enable_variable_to_check_98[5] = enable_variable_233_to_check_98;


// 校验节点99的接口
wire [35:0] value_variable_to_check_99;
wire [35:0] value_check_99_to_variable;
wire [5:0] enable_variable_to_check_99;
wire [5:0] enable_check_99_to_variable;

// 拆分后校验节点99传递给变量节点2的值以及对变量节点2传递过来的值
wire [5:0] value_check_99_to_variable_2;
wire enable_check_99_to_variable_2;
wire [5:0] value_variable_2_to_check_99;
wire enable_variable_2_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_2 = value_check_99_to_variable[5:0];
assign enable_check_99_to_variable_2 = enable_check_99_to_variable[0];
// 对变量节点2传递过来的值进行组合
assign value_variable_to_check_99[5:0] = value_variable_2_to_check_99;
assign enable_variable_to_check_99[0] = enable_variable_2_to_check_99;

// 拆分后校验节点99传递给变量节点83的值以及对变量节点83传递过来的值
wire [5:0] value_check_99_to_variable_83;
wire enable_check_99_to_variable_83;
wire [5:0] value_variable_83_to_check_99;
wire enable_variable_83_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_83 = value_check_99_to_variable[11:6];
assign enable_check_99_to_variable_83 = enable_check_99_to_variable[1];
// 对变量节点83传递过来的值进行组合
assign value_variable_to_check_99[11:6] = value_variable_83_to_check_99;
assign enable_variable_to_check_99[1] = enable_variable_83_to_check_99;

// 拆分后校验节点99传递给变量节点117的值以及对变量节点117传递过来的值
wire [5:0] value_check_99_to_variable_117;
wire enable_check_99_to_variable_117;
wire [5:0] value_variable_117_to_check_99;
wire enable_variable_117_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_117 = value_check_99_to_variable[17:12];
assign enable_check_99_to_variable_117 = enable_check_99_to_variable[2];
// 对变量节点117传递过来的值进行组合
assign value_variable_to_check_99[17:12] = value_variable_117_to_check_99;
assign enable_variable_to_check_99[2] = enable_variable_117_to_check_99;

// 拆分后校验节点99传递给变量节点168的值以及对变量节点168传递过来的值
wire [5:0] value_check_99_to_variable_168;
wire enable_check_99_to_variable_168;
wire [5:0] value_variable_168_to_check_99;
wire enable_variable_168_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_168 = value_check_99_to_variable[23:18];
assign enable_check_99_to_variable_168 = enable_check_99_to_variable[3];
// 对变量节点168传递过来的值进行组合
assign value_variable_to_check_99[23:18] = value_variable_168_to_check_99;
assign enable_variable_to_check_99[3] = enable_variable_168_to_check_99;

// 拆分后校验节点99传递给变量节点212的值以及对变量节点212传递过来的值
wire [5:0] value_check_99_to_variable_212;
wire enable_check_99_to_variable_212;
wire [5:0] value_variable_212_to_check_99;
wire enable_variable_212_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_212 = value_check_99_to_variable[29:24];
assign enable_check_99_to_variable_212 = enable_check_99_to_variable[4];
// 对变量节点212传递过来的值进行组合
assign value_variable_to_check_99[29:24] = value_variable_212_to_check_99;
assign enable_variable_to_check_99[4] = enable_variable_212_to_check_99;

// 拆分后校验节点99传递给变量节点215的值以及对变量节点215传递过来的值
wire [5:0] value_check_99_to_variable_215;
wire enable_check_99_to_variable_215;
wire [5:0] value_variable_215_to_check_99;
wire enable_variable_215_to_check_99;
// 对校验节点99的输出值进行拆分
assign value_check_99_to_variable_215 = value_check_99_to_variable[35:30];
assign enable_check_99_to_variable_215 = enable_check_99_to_variable[5];
// 对变量节点215传递过来的值进行组合
assign value_variable_to_check_99[35:30] = value_variable_215_to_check_99;
assign enable_variable_to_check_99[5] = enable_variable_215_to_check_99;


// 校验节点100的接口
wire [35:0] value_variable_to_check_100;
wire [35:0] value_check_100_to_variable;
wire [5:0] enable_variable_to_check_100;
wire [5:0] enable_check_100_to_variable;

// 拆分后校验节点100传递给变量节点0的值以及对变量节点0传递过来的值
wire [5:0] value_check_100_to_variable_0;
wire enable_check_100_to_variable_0;
wire [5:0] value_variable_0_to_check_100;
wire enable_variable_0_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_0 = value_check_100_to_variable[5:0];
assign enable_check_100_to_variable_0 = enable_check_100_to_variable[0];
// 对变量节点0传递过来的值进行组合
assign value_variable_to_check_100[5:0] = value_variable_0_to_check_100;
assign enable_variable_to_check_100[0] = enable_variable_0_to_check_100;

// 拆分后校验节点100传递给变量节点84的值以及对变量节点84传递过来的值
wire [5:0] value_check_100_to_variable_84;
wire enable_check_100_to_variable_84;
wire [5:0] value_variable_84_to_check_100;
wire enable_variable_84_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_84 = value_check_100_to_variable[11:6];
assign enable_check_100_to_variable_84 = enable_check_100_to_variable[1];
// 对变量节点84传递过来的值进行组合
assign value_variable_to_check_100[11:6] = value_variable_84_to_check_100;
assign enable_variable_to_check_100[1] = enable_variable_84_to_check_100;

// 拆分后校验节点100传递给变量节点115的值以及对变量节点115传递过来的值
wire [5:0] value_check_100_to_variable_115;
wire enable_check_100_to_variable_115;
wire [5:0] value_variable_115_to_check_100;
wire enable_variable_115_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_115 = value_check_100_to_variable[17:12];
assign enable_check_100_to_variable_115 = enable_check_100_to_variable[2];
// 对变量节点115传递过来的值进行组合
assign value_variable_to_check_100[17:12] = value_variable_115_to_check_100;
assign enable_variable_to_check_100[2] = enable_variable_115_to_check_100;

// 拆分后校验节点100传递给变量节点166的值以及对变量节点166传递过来的值
wire [5:0] value_check_100_to_variable_166;
wire enable_check_100_to_variable_166;
wire [5:0] value_variable_166_to_check_100;
wire enable_variable_166_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_166 = value_check_100_to_variable[23:18];
assign enable_check_100_to_variable_166 = enable_check_100_to_variable[3];
// 对变量节点166传递过来的值进行组合
assign value_variable_to_check_100[23:18] = value_variable_166_to_check_100;
assign enable_variable_to_check_100[3] = enable_variable_166_to_check_100;

// 拆分后校验节点100传递给变量节点203的值以及对变量节点203传递过来的值
wire [5:0] value_check_100_to_variable_203;
wire enable_check_100_to_variable_203;
wire [5:0] value_variable_203_to_check_100;
wire enable_variable_203_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_203 = value_check_100_to_variable[29:24];
assign enable_check_100_to_variable_203 = enable_check_100_to_variable[4];
// 对变量节点203传递过来的值进行组合
assign value_variable_to_check_100[29:24] = value_variable_203_to_check_100;
assign enable_variable_to_check_100[4] = enable_variable_203_to_check_100;

// 拆分后校验节点100传递给变量节点223的值以及对变量节点223传递过来的值
wire [5:0] value_check_100_to_variable_223;
wire enable_check_100_to_variable_223;
wire [5:0] value_variable_223_to_check_100;
wire enable_variable_223_to_check_100;
// 对校验节点100的输出值进行拆分
assign value_check_100_to_variable_223 = value_check_100_to_variable[35:30];
assign enable_check_100_to_variable_223 = enable_check_100_to_variable[5];
// 对变量节点223传递过来的值进行组合
assign value_variable_to_check_100[35:30] = value_variable_223_to_check_100;
assign enable_variable_to_check_100[5] = enable_variable_223_to_check_100;


// 校验节点101的接口
wire [35:0] value_variable_to_check_101;
wire [35:0] value_check_101_to_variable;
wire [5:0] enable_variable_to_check_101;
wire [5:0] enable_check_101_to_variable;

// 拆分后校验节点101传递给变量节点4的值以及对变量节点4传递过来的值
wire [5:0] value_check_101_to_variable_4;
wire enable_check_101_to_variable_4;
wire [5:0] value_variable_4_to_check_101;
wire enable_variable_4_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_4 = value_check_101_to_variable[5:0];
assign enable_check_101_to_variable_4 = enable_check_101_to_variable[0];
// 对变量节点4传递过来的值进行组合
assign value_variable_to_check_101[5:0] = value_variable_4_to_check_101;
assign enable_variable_to_check_101[0] = enable_variable_4_to_check_101;

// 拆分后校验节点101传递给变量节点80的值以及对变量节点80传递过来的值
wire [5:0] value_check_101_to_variable_80;
wire enable_check_101_to_variable_80;
wire [5:0] value_variable_80_to_check_101;
wire enable_variable_80_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_80 = value_check_101_to_variable[11:6];
assign enable_check_101_to_variable_80 = enable_check_101_to_variable[1];
// 对变量节点80传递过来的值进行组合
assign value_variable_to_check_101[11:6] = value_variable_80_to_check_101;
assign enable_variable_to_check_101[1] = enable_variable_80_to_check_101;

// 拆分后校验节点101传递给变量节点99的值以及对变量节点99传递过来的值
wire [5:0] value_check_101_to_variable_99;
wire enable_check_101_to_variable_99;
wire [5:0] value_variable_99_to_check_101;
wire enable_variable_99_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_99 = value_check_101_to_variable[17:12];
assign enable_check_101_to_variable_99 = enable_check_101_to_variable[2];
// 对变量节点99传递过来的值进行组合
assign value_variable_to_check_101[17:12] = value_variable_99_to_check_101;
assign enable_variable_to_check_101[2] = enable_variable_99_to_check_101;

// 拆分后校验节点101传递给变量节点158的值以及对变量节点158传递过来的值
wire [5:0] value_check_101_to_variable_158;
wire enable_check_101_to_variable_158;
wire [5:0] value_variable_158_to_check_101;
wire enable_variable_158_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_158 = value_check_101_to_variable[23:18];
assign enable_check_101_to_variable_158 = enable_check_101_to_variable[3];
// 对变量节点158传递过来的值进行组合
assign value_variable_to_check_101[23:18] = value_variable_158_to_check_101;
assign enable_variable_to_check_101[3] = enable_variable_158_to_check_101;

// 拆分后校验节点101传递给变量节点181的值以及对变量节点181传递过来的值
wire [5:0] value_check_101_to_variable_181;
wire enable_check_101_to_variable_181;
wire [5:0] value_variable_181_to_check_101;
wire enable_variable_181_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_181 = value_check_101_to_variable[29:24];
assign enable_check_101_to_variable_181 = enable_check_101_to_variable[4];
// 对变量节点181传递过来的值进行组合
assign value_variable_to_check_101[29:24] = value_variable_181_to_check_101;
assign enable_variable_to_check_101[4] = enable_variable_181_to_check_101;

// 拆分后校验节点101传递给变量节点221的值以及对变量节点221传递过来的值
wire [5:0] value_check_101_to_variable_221;
wire enable_check_101_to_variable_221;
wire [5:0] value_variable_221_to_check_101;
wire enable_variable_221_to_check_101;
// 对校验节点101的输出值进行拆分
assign value_check_101_to_variable_221 = value_check_101_to_variable[35:30];
assign enable_check_101_to_variable_221 = enable_check_101_to_variable[5];
// 对变量节点221传递过来的值进行组合
assign value_variable_to_check_101[35:30] = value_variable_221_to_check_101;
assign enable_variable_to_check_101[5] = enable_variable_221_to_check_101;


// 校验节点102的接口
wire [35:0] value_variable_to_check_102;
wire [35:0] value_check_102_to_variable;
wire [5:0] enable_variable_to_check_102;
wire [5:0] enable_check_102_to_variable;

// 拆分后校验节点102传递给变量节点41的值以及对变量节点41传递过来的值
wire [5:0] value_check_102_to_variable_41;
wire enable_check_102_to_variable_41;
wire [5:0] value_variable_41_to_check_102;
wire enable_variable_41_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_41 = value_check_102_to_variable[5:0];
assign enable_check_102_to_variable_41 = enable_check_102_to_variable[0];
// 对变量节点41传递过来的值进行组合
assign value_variable_to_check_102[5:0] = value_variable_41_to_check_102;
assign enable_variable_to_check_102[0] = enable_variable_41_to_check_102;

// 拆分后校验节点102传递给变量节点68的值以及对变量节点68传递过来的值
wire [5:0] value_check_102_to_variable_68;
wire enable_check_102_to_variable_68;
wire [5:0] value_variable_68_to_check_102;
wire enable_variable_68_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_68 = value_check_102_to_variable[11:6];
assign enable_check_102_to_variable_68 = enable_check_102_to_variable[1];
// 对变量节点68传递过来的值进行组合
assign value_variable_to_check_102[11:6] = value_variable_68_to_check_102;
assign enable_variable_to_check_102[1] = enable_variable_68_to_check_102;

// 拆分后校验节点102传递给变量节点115的值以及对变量节点115传递过来的值
wire [5:0] value_check_102_to_variable_115;
wire enable_check_102_to_variable_115;
wire [5:0] value_variable_115_to_check_102;
wire enable_variable_115_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_115 = value_check_102_to_variable[17:12];
assign enable_check_102_to_variable_115 = enable_check_102_to_variable[2];
// 对变量节点115传递过来的值进行组合
assign value_variable_to_check_102[17:12] = value_variable_115_to_check_102;
assign enable_variable_to_check_102[2] = enable_variable_115_to_check_102;

// 拆分后校验节点102传递给变量节点148的值以及对变量节点148传递过来的值
wire [5:0] value_check_102_to_variable_148;
wire enable_check_102_to_variable_148;
wire [5:0] value_variable_148_to_check_102;
wire enable_variable_148_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_148 = value_check_102_to_variable[23:18];
assign enable_check_102_to_variable_148 = enable_check_102_to_variable[3];
// 对变量节点148传递过来的值进行组合
assign value_variable_to_check_102[23:18] = value_variable_148_to_check_102;
assign enable_variable_to_check_102[3] = enable_variable_148_to_check_102;

// 拆分后校验节点102传递给变量节点196的值以及对变量节点196传递过来的值
wire [5:0] value_check_102_to_variable_196;
wire enable_check_102_to_variable_196;
wire [5:0] value_variable_196_to_check_102;
wire enable_variable_196_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_196 = value_check_102_to_variable[29:24];
assign enable_check_102_to_variable_196 = enable_check_102_to_variable[4];
// 对变量节点196传递过来的值进行组合
assign value_variable_to_check_102[29:24] = value_variable_196_to_check_102;
assign enable_variable_to_check_102[4] = enable_variable_196_to_check_102;

// 拆分后校验节点102传递给变量节点229的值以及对变量节点229传递过来的值
wire [5:0] value_check_102_to_variable_229;
wire enable_check_102_to_variable_229;
wire [5:0] value_variable_229_to_check_102;
wire enable_variable_229_to_check_102;
// 对校验节点102的输出值进行拆分
assign value_check_102_to_variable_229 = value_check_102_to_variable[35:30];
assign enable_check_102_to_variable_229 = enable_check_102_to_variable[5];
// 对变量节点229传递过来的值进行组合
assign value_variable_to_check_102[35:30] = value_variable_229_to_check_102;
assign enable_variable_to_check_102[5] = enable_variable_229_to_check_102;


// 校验节点103的接口
wire [35:0] value_variable_to_check_103;
wire [35:0] value_check_103_to_variable;
wire [5:0] enable_variable_to_check_103;
wire [5:0] enable_check_103_to_variable;

// 拆分后校验节点103传递给变量节点38的值以及对变量节点38传递过来的值
wire [5:0] value_check_103_to_variable_38;
wire enable_check_103_to_variable_38;
wire [5:0] value_variable_38_to_check_103;
wire enable_variable_38_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_38 = value_check_103_to_variable[5:0];
assign enable_check_103_to_variable_38 = enable_check_103_to_variable[0];
// 对变量节点38传递过来的值进行组合
assign value_variable_to_check_103[5:0] = value_variable_38_to_check_103;
assign enable_variable_to_check_103[0] = enable_variable_38_to_check_103;

// 拆分后校验节点103传递给变量节点73的值以及对变量节点73传递过来的值
wire [5:0] value_check_103_to_variable_73;
wire enable_check_103_to_variable_73;
wire [5:0] value_variable_73_to_check_103;
wire enable_variable_73_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_73 = value_check_103_to_variable[11:6];
assign enable_check_103_to_variable_73 = enable_check_103_to_variable[1];
// 对变量节点73传递过来的值进行组合
assign value_variable_to_check_103[11:6] = value_variable_73_to_check_103;
assign enable_variable_to_check_103[1] = enable_variable_73_to_check_103;

// 拆分后校验节点103传递给变量节点102的值以及对变量节点102传递过来的值
wire [5:0] value_check_103_to_variable_102;
wire enable_check_103_to_variable_102;
wire [5:0] value_variable_102_to_check_103;
wire enable_variable_102_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_102 = value_check_103_to_variable[17:12];
assign enable_check_103_to_variable_102 = enable_check_103_to_variable[2];
// 对变量节点102传递过来的值进行组合
assign value_variable_to_check_103[17:12] = value_variable_102_to_check_103;
assign enable_variable_to_check_103[2] = enable_variable_102_to_check_103;

// 拆分后校验节点103传递给变量节点165的值以及对变量节点165传递过来的值
wire [5:0] value_check_103_to_variable_165;
wire enable_check_103_to_variable_165;
wire [5:0] value_variable_165_to_check_103;
wire enable_variable_165_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_165 = value_check_103_to_variable[23:18];
assign enable_check_103_to_variable_165 = enable_check_103_to_variable[3];
// 对变量节点165传递过来的值进行组合
assign value_variable_to_check_103[23:18] = value_variable_165_to_check_103;
assign enable_variable_to_check_103[3] = enable_variable_165_to_check_103;

// 拆分后校验节点103传递给变量节点192的值以及对变量节点192传递过来的值
wire [5:0] value_check_103_to_variable_192;
wire enable_check_103_to_variable_192;
wire [5:0] value_variable_192_to_check_103;
wire enable_variable_192_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_192 = value_check_103_to_variable[29:24];
assign enable_check_103_to_variable_192 = enable_check_103_to_variable[4];
// 对变量节点192传递过来的值进行组合
assign value_variable_to_check_103[29:24] = value_variable_192_to_check_103;
assign enable_variable_to_check_103[4] = enable_variable_192_to_check_103;

// 拆分后校验节点103传递给变量节点251的值以及对变量节点251传递过来的值
wire [5:0] value_check_103_to_variable_251;
wire enable_check_103_to_variable_251;
wire [5:0] value_variable_251_to_check_103;
wire enable_variable_251_to_check_103;
// 对校验节点103的输出值进行拆分
assign value_check_103_to_variable_251 = value_check_103_to_variable[35:30];
assign enable_check_103_to_variable_251 = enable_check_103_to_variable[5];
// 对变量节点251传递过来的值进行组合
assign value_variable_to_check_103[35:30] = value_variable_251_to_check_103;
assign enable_variable_to_check_103[5] = enable_variable_251_to_check_103;


// 校验节点104的接口
wire [35:0] value_variable_to_check_104;
wire [35:0] value_check_104_to_variable;
wire [5:0] enable_variable_to_check_104;
wire [5:0] enable_check_104_to_variable;

// 拆分后校验节点104传递给变量节点17的值以及对变量节点17传递过来的值
wire [5:0] value_check_104_to_variable_17;
wire enable_check_104_to_variable_17;
wire [5:0] value_variable_17_to_check_104;
wire enable_variable_17_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_17 = value_check_104_to_variable[5:0];
assign enable_check_104_to_variable_17 = enable_check_104_to_variable[0];
// 对变量节点17传递过来的值进行组合
assign value_variable_to_check_104[5:0] = value_variable_17_to_check_104;
assign enable_variable_to_check_104[0] = enable_variable_17_to_check_104;

// 拆分后校验节点104传递给变量节点83的值以及对变量节点83传递过来的值
wire [5:0] value_check_104_to_variable_83;
wire enable_check_104_to_variable_83;
wire [5:0] value_variable_83_to_check_104;
wire enable_variable_83_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_83 = value_check_104_to_variable[11:6];
assign enable_check_104_to_variable_83 = enable_check_104_to_variable[1];
// 对变量节点83传递过来的值进行组合
assign value_variable_to_check_104[11:6] = value_variable_83_to_check_104;
assign enable_variable_to_check_104[1] = enable_variable_83_to_check_104;

// 拆分后校验节点104传递给变量节点123的值以及对变量节点123传递过来的值
wire [5:0] value_check_104_to_variable_123;
wire enable_check_104_to_variable_123;
wire [5:0] value_variable_123_to_check_104;
wire enable_variable_123_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_123 = value_check_104_to_variable[17:12];
assign enable_check_104_to_variable_123 = enable_check_104_to_variable[2];
// 对变量节点123传递过来的值进行组合
assign value_variable_to_check_104[17:12] = value_variable_123_to_check_104;
assign enable_variable_to_check_104[2] = enable_variable_123_to_check_104;

// 拆分后校验节点104传递给变量节点144的值以及对变量节点144传递过来的值
wire [5:0] value_check_104_to_variable_144;
wire enable_check_104_to_variable_144;
wire [5:0] value_variable_144_to_check_104;
wire enable_variable_144_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_144 = value_check_104_to_variable[23:18];
assign enable_check_104_to_variable_144 = enable_check_104_to_variable[3];
// 对变量节点144传递过来的值进行组合
assign value_variable_to_check_104[23:18] = value_variable_144_to_check_104;
assign enable_variable_to_check_104[3] = enable_variable_144_to_check_104;

// 拆分后校验节点104传递给变量节点205的值以及对变量节点205传递过来的值
wire [5:0] value_check_104_to_variable_205;
wire enable_check_104_to_variable_205;
wire [5:0] value_variable_205_to_check_104;
wire enable_variable_205_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_205 = value_check_104_to_variable[29:24];
assign enable_check_104_to_variable_205 = enable_check_104_to_variable[4];
// 对变量节点205传递过来的值进行组合
assign value_variable_to_check_104[29:24] = value_variable_205_to_check_104;
assign enable_variable_to_check_104[4] = enable_variable_205_to_check_104;

// 拆分后校验节点104传递给变量节点237的值以及对变量节点237传递过来的值
wire [5:0] value_check_104_to_variable_237;
wire enable_check_104_to_variable_237;
wire [5:0] value_variable_237_to_check_104;
wire enable_variable_237_to_check_104;
// 对校验节点104的输出值进行拆分
assign value_check_104_to_variable_237 = value_check_104_to_variable[35:30];
assign enable_check_104_to_variable_237 = enable_check_104_to_variable[5];
// 对变量节点237传递过来的值进行组合
assign value_variable_to_check_104[35:30] = value_variable_237_to_check_104;
assign enable_variable_to_check_104[5] = enable_variable_237_to_check_104;


// 校验节点105的接口
wire [35:0] value_variable_to_check_105;
wire [35:0] value_check_105_to_variable;
wire [5:0] enable_variable_to_check_105;
wire [5:0] enable_check_105_to_variable;

// 拆分后校验节点105传递给变量节点19的值以及对变量节点19传递过来的值
wire [5:0] value_check_105_to_variable_19;
wire enable_check_105_to_variable_19;
wire [5:0] value_variable_19_to_check_105;
wire enable_variable_19_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_19 = value_check_105_to_variable[5:0];
assign enable_check_105_to_variable_19 = enable_check_105_to_variable[0];
// 对变量节点19传递过来的值进行组合
assign value_variable_to_check_105[5:0] = value_variable_19_to_check_105;
assign enable_variable_to_check_105[0] = enable_variable_19_to_check_105;

// 拆分后校验节点105传递给变量节点83的值以及对变量节点83传递过来的值
wire [5:0] value_check_105_to_variable_83;
wire enable_check_105_to_variable_83;
wire [5:0] value_variable_83_to_check_105;
wire enable_variable_83_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_83 = value_check_105_to_variable[11:6];
assign enable_check_105_to_variable_83 = enable_check_105_to_variable[1];
// 对变量节点83传递过来的值进行组合
assign value_variable_to_check_105[11:6] = value_variable_83_to_check_105;
assign enable_variable_to_check_105[1] = enable_variable_83_to_check_105;

// 拆分后校验节点105传递给变量节点93的值以及对变量节点93传递过来的值
wire [5:0] value_check_105_to_variable_93;
wire enable_check_105_to_variable_93;
wire [5:0] value_variable_93_to_check_105;
wire enable_variable_93_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_93 = value_check_105_to_variable[17:12];
assign enable_check_105_to_variable_93 = enable_check_105_to_variable[2];
// 对变量节点93传递过来的值进行组合
assign value_variable_to_check_105[17:12] = value_variable_93_to_check_105;
assign enable_variable_to_check_105[2] = enable_variable_93_to_check_105;

// 拆分后校验节点105传递给变量节点170的值以及对变量节点170传递过来的值
wire [5:0] value_check_105_to_variable_170;
wire enable_check_105_to_variable_170;
wire [5:0] value_variable_170_to_check_105;
wire enable_variable_170_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_170 = value_check_105_to_variable[23:18];
assign enable_check_105_to_variable_170 = enable_check_105_to_variable[3];
// 对变量节点170传递过来的值进行组合
assign value_variable_to_check_105[23:18] = value_variable_170_to_check_105;
assign enable_variable_to_check_105[3] = enable_variable_170_to_check_105;

// 拆分后校验节点105传递给变量节点204的值以及对变量节点204传递过来的值
wire [5:0] value_check_105_to_variable_204;
wire enable_check_105_to_variable_204;
wire [5:0] value_variable_204_to_check_105;
wire enable_variable_204_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_204 = value_check_105_to_variable[29:24];
assign enable_check_105_to_variable_204 = enable_check_105_to_variable[4];
// 对变量节点204传递过来的值进行组合
assign value_variable_to_check_105[29:24] = value_variable_204_to_check_105;
assign enable_variable_to_check_105[4] = enable_variable_204_to_check_105;

// 拆分后校验节点105传递给变量节点249的值以及对变量节点249传递过来的值
wire [5:0] value_check_105_to_variable_249;
wire enable_check_105_to_variable_249;
wire [5:0] value_variable_249_to_check_105;
wire enable_variable_249_to_check_105;
// 对校验节点105的输出值进行拆分
assign value_check_105_to_variable_249 = value_check_105_to_variable[35:30];
assign enable_check_105_to_variable_249 = enable_check_105_to_variable[5];
// 对变量节点249传递过来的值进行组合
assign value_variable_to_check_105[35:30] = value_variable_249_to_check_105;
assign enable_variable_to_check_105[5] = enable_variable_249_to_check_105;


// 校验节点106的接口
wire [35:0] value_variable_to_check_106;
wire [35:0] value_check_106_to_variable;
wire [5:0] enable_variable_to_check_106;
wire [5:0] enable_check_106_to_variable;

// 拆分后校验节点106传递给变量节点1的值以及对变量节点1传递过来的值
wire [5:0] value_check_106_to_variable_1;
wire enable_check_106_to_variable_1;
wire [5:0] value_variable_1_to_check_106;
wire enable_variable_1_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_1 = value_check_106_to_variable[5:0];
assign enable_check_106_to_variable_1 = enable_check_106_to_variable[0];
// 对变量节点1传递过来的值进行组合
assign value_variable_to_check_106[5:0] = value_variable_1_to_check_106;
assign enable_variable_to_check_106[0] = enable_variable_1_to_check_106;

// 拆分后校验节点106传递给变量节点75的值以及对变量节点75传递过来的值
wire [5:0] value_check_106_to_variable_75;
wire enable_check_106_to_variable_75;
wire [5:0] value_variable_75_to_check_106;
wire enable_variable_75_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_75 = value_check_106_to_variable[11:6];
assign enable_check_106_to_variable_75 = enable_check_106_to_variable[1];
// 对变量节点75传递过来的值进行组合
assign value_variable_to_check_106[11:6] = value_variable_75_to_check_106;
assign enable_variable_to_check_106[1] = enable_variable_75_to_check_106;

// 拆分后校验节点106传递给变量节点127的值以及对变量节点127传递过来的值
wire [5:0] value_check_106_to_variable_127;
wire enable_check_106_to_variable_127;
wire [5:0] value_variable_127_to_check_106;
wire enable_variable_127_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_127 = value_check_106_to_variable[17:12];
assign enable_check_106_to_variable_127 = enable_check_106_to_variable[2];
// 对变量节点127传递过来的值进行组合
assign value_variable_to_check_106[17:12] = value_variable_127_to_check_106;
assign enable_variable_to_check_106[2] = enable_variable_127_to_check_106;

// 拆分后校验节点106传递给变量节点166的值以及对变量节点166传递过来的值
wire [5:0] value_check_106_to_variable_166;
wire enable_check_106_to_variable_166;
wire [5:0] value_variable_166_to_check_106;
wire enable_variable_166_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_166 = value_check_106_to_variable[23:18];
assign enable_check_106_to_variable_166 = enable_check_106_to_variable[3];
// 对变量节点166传递过来的值进行组合
assign value_variable_to_check_106[23:18] = value_variable_166_to_check_106;
assign enable_variable_to_check_106[3] = enable_variable_166_to_check_106;

// 拆分后校验节点106传递给变量节点200的值以及对变量节点200传递过来的值
wire [5:0] value_check_106_to_variable_200;
wire enable_check_106_to_variable_200;
wire [5:0] value_variable_200_to_check_106;
wire enable_variable_200_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_200 = value_check_106_to_variable[29:24];
assign enable_check_106_to_variable_200 = enable_check_106_to_variable[4];
// 对变量节点200传递过来的值进行组合
assign value_variable_to_check_106[29:24] = value_variable_200_to_check_106;
assign enable_variable_to_check_106[4] = enable_variable_200_to_check_106;

// 拆分后校验节点106传递给变量节点254的值以及对变量节点254传递过来的值
wire [5:0] value_check_106_to_variable_254;
wire enable_check_106_to_variable_254;
wire [5:0] value_variable_254_to_check_106;
wire enable_variable_254_to_check_106;
// 对校验节点106的输出值进行拆分
assign value_check_106_to_variable_254 = value_check_106_to_variable[35:30];
assign enable_check_106_to_variable_254 = enable_check_106_to_variable[5];
// 对变量节点254传递过来的值进行组合
assign value_variable_to_check_106[35:30] = value_variable_254_to_check_106;
assign enable_variable_to_check_106[5] = enable_variable_254_to_check_106;


// 校验节点107的接口
wire [35:0] value_variable_to_check_107;
wire [35:0] value_check_107_to_variable;
wire [5:0] enable_variable_to_check_107;
wire [5:0] enable_check_107_to_variable;

// 拆分后校验节点107传递给变量节点10的值以及对变量节点10传递过来的值
wire [5:0] value_check_107_to_variable_10;
wire enable_check_107_to_variable_10;
wire [5:0] value_variable_10_to_check_107;
wire enable_variable_10_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_10 = value_check_107_to_variable[5:0];
assign enable_check_107_to_variable_10 = enable_check_107_to_variable[0];
// 对变量节点10传递过来的值进行组合
assign value_variable_to_check_107[5:0] = value_variable_10_to_check_107;
assign enable_variable_to_check_107[0] = enable_variable_10_to_check_107;

// 拆分后校验节点107传递给变量节点54的值以及对变量节点54传递过来的值
wire [5:0] value_check_107_to_variable_54;
wire enable_check_107_to_variable_54;
wire [5:0] value_variable_54_to_check_107;
wire enable_variable_54_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_54 = value_check_107_to_variable[11:6];
assign enable_check_107_to_variable_54 = enable_check_107_to_variable[1];
// 对变量节点54传递过来的值进行组合
assign value_variable_to_check_107[11:6] = value_variable_54_to_check_107;
assign enable_variable_to_check_107[1] = enable_variable_54_to_check_107;

// 拆分后校验节点107传递给变量节点118的值以及对变量节点118传递过来的值
wire [5:0] value_check_107_to_variable_118;
wire enable_check_107_to_variable_118;
wire [5:0] value_variable_118_to_check_107;
wire enable_variable_118_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_118 = value_check_107_to_variable[17:12];
assign enable_check_107_to_variable_118 = enable_check_107_to_variable[2];
// 对变量节点118传递过来的值进行组合
assign value_variable_to_check_107[17:12] = value_variable_118_to_check_107;
assign enable_variable_to_check_107[2] = enable_variable_118_to_check_107;

// 拆分后校验节点107传递给变量节点162的值以及对变量节点162传递过来的值
wire [5:0] value_check_107_to_variable_162;
wire enable_check_107_to_variable_162;
wire [5:0] value_variable_162_to_check_107;
wire enable_variable_162_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_162 = value_check_107_to_variable[23:18];
assign enable_check_107_to_variable_162 = enable_check_107_to_variable[3];
// 对变量节点162传递过来的值进行组合
assign value_variable_to_check_107[23:18] = value_variable_162_to_check_107;
assign enable_variable_to_check_107[3] = enable_variable_162_to_check_107;

// 拆分后校验节点107传递给变量节点213的值以及对变量节点213传递过来的值
wire [5:0] value_check_107_to_variable_213;
wire enable_check_107_to_variable_213;
wire [5:0] value_variable_213_to_check_107;
wire enable_variable_213_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_213 = value_check_107_to_variable[29:24];
assign enable_check_107_to_variable_213 = enable_check_107_to_variable[4];
// 对变量节点213传递过来的值进行组合
assign value_variable_to_check_107[29:24] = value_variable_213_to_check_107;
assign enable_variable_to_check_107[4] = enable_variable_213_to_check_107;

// 拆分后校验节点107传递给变量节点222的值以及对变量节点222传递过来的值
wire [5:0] value_check_107_to_variable_222;
wire enable_check_107_to_variable_222;
wire [5:0] value_variable_222_to_check_107;
wire enable_variable_222_to_check_107;
// 对校验节点107的输出值进行拆分
assign value_check_107_to_variable_222 = value_check_107_to_variable[35:30];
assign enable_check_107_to_variable_222 = enable_check_107_to_variable[5];
// 对变量节点222传递过来的值进行组合
assign value_variable_to_check_107[35:30] = value_variable_222_to_check_107;
assign enable_variable_to_check_107[5] = enable_variable_222_to_check_107;


// 校验节点108的接口
wire [35:0] value_variable_to_check_108;
wire [35:0] value_check_108_to_variable;
wire [5:0] enable_variable_to_check_108;
wire [5:0] enable_check_108_to_variable;

// 拆分后校验节点108传递给变量节点40的值以及对变量节点40传递过来的值
wire [5:0] value_check_108_to_variable_40;
wire enable_check_108_to_variable_40;
wire [5:0] value_variable_40_to_check_108;
wire enable_variable_40_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_40 = value_check_108_to_variable[5:0];
assign enable_check_108_to_variable_40 = enable_check_108_to_variable[0];
// 对变量节点40传递过来的值进行组合
assign value_variable_to_check_108[5:0] = value_variable_40_to_check_108;
assign enable_variable_to_check_108[0] = enable_variable_40_to_check_108;

// 拆分后校验节点108传递给变量节点81的值以及对变量节点81传递过来的值
wire [5:0] value_check_108_to_variable_81;
wire enable_check_108_to_variable_81;
wire [5:0] value_variable_81_to_check_108;
wire enable_variable_81_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_81 = value_check_108_to_variable[11:6];
assign enable_check_108_to_variable_81 = enable_check_108_to_variable[1];
// 对变量节点81传递过来的值进行组合
assign value_variable_to_check_108[11:6] = value_variable_81_to_check_108;
assign enable_variable_to_check_108[1] = enable_variable_81_to_check_108;

// 拆分后校验节点108传递给变量节点126的值以及对变量节点126传递过来的值
wire [5:0] value_check_108_to_variable_126;
wire enable_check_108_to_variable_126;
wire [5:0] value_variable_126_to_check_108;
wire enable_variable_126_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_126 = value_check_108_to_variable[17:12];
assign enable_check_108_to_variable_126 = enable_check_108_to_variable[2];
// 对变量节点126传递过来的值进行组合
assign value_variable_to_check_108[17:12] = value_variable_126_to_check_108;
assign enable_variable_to_check_108[2] = enable_variable_126_to_check_108;

// 拆分后校验节点108传递给变量节点169的值以及对变量节点169传递过来的值
wire [5:0] value_check_108_to_variable_169;
wire enable_check_108_to_variable_169;
wire [5:0] value_variable_169_to_check_108;
wire enable_variable_169_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_169 = value_check_108_to_variable[23:18];
assign enable_check_108_to_variable_169 = enable_check_108_to_variable[3];
// 对变量节点169传递过来的值进行组合
assign value_variable_to_check_108[23:18] = value_variable_169_to_check_108;
assign enable_variable_to_check_108[3] = enable_variable_169_to_check_108;

// 拆分后校验节点108传递给变量节点210的值以及对变量节点210传递过来的值
wire [5:0] value_check_108_to_variable_210;
wire enable_check_108_to_variable_210;
wire [5:0] value_variable_210_to_check_108;
wire enable_variable_210_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_210 = value_check_108_to_variable[29:24];
assign enable_check_108_to_variable_210 = enable_check_108_to_variable[4];
// 对变量节点210传递过来的值进行组合
assign value_variable_to_check_108[29:24] = value_variable_210_to_check_108;
assign enable_variable_to_check_108[4] = enable_variable_210_to_check_108;

// 拆分后校验节点108传递给变量节点253的值以及对变量节点253传递过来的值
wire [5:0] value_check_108_to_variable_253;
wire enable_check_108_to_variable_253;
wire [5:0] value_variable_253_to_check_108;
wire enable_variable_253_to_check_108;
// 对校验节点108的输出值进行拆分
assign value_check_108_to_variable_253 = value_check_108_to_variable[35:30];
assign enable_check_108_to_variable_253 = enable_check_108_to_variable[5];
// 对变量节点253传递过来的值进行组合
assign value_variable_to_check_108[35:30] = value_variable_253_to_check_108;
assign enable_variable_to_check_108[5] = enable_variable_253_to_check_108;


// 校验节点109的接口
wire [35:0] value_variable_to_check_109;
wire [35:0] value_check_109_to_variable;
wire [5:0] enable_variable_to_check_109;
wire [5:0] enable_check_109_to_variable;

// 拆分后校验节点109传递给变量节点34的值以及对变量节点34传递过来的值
wire [5:0] value_check_109_to_variable_34;
wire enable_check_109_to_variable_34;
wire [5:0] value_variable_34_to_check_109;
wire enable_variable_34_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_34 = value_check_109_to_variable[5:0];
assign enable_check_109_to_variable_34 = enable_check_109_to_variable[0];
// 对变量节点34传递过来的值进行组合
assign value_variable_to_check_109[5:0] = value_variable_34_to_check_109;
assign enable_variable_to_check_109[0] = enable_variable_34_to_check_109;

// 拆分后校验节点109传递给变量节点85的值以及对变量节点85传递过来的值
wire [5:0] value_check_109_to_variable_85;
wire enable_check_109_to_variable_85;
wire [5:0] value_variable_85_to_check_109;
wire enable_variable_85_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_85 = value_check_109_to_variable[11:6];
assign enable_check_109_to_variable_85 = enable_check_109_to_variable[1];
// 对变量节点85传递过来的值进行组合
assign value_variable_to_check_109[11:6] = value_variable_85_to_check_109;
assign enable_variable_to_check_109[1] = enable_variable_85_to_check_109;

// 拆分后校验节点109传递给变量节点116的值以及对变量节点116传递过来的值
wire [5:0] value_check_109_to_variable_116;
wire enable_check_109_to_variable_116;
wire [5:0] value_variable_116_to_check_109;
wire enable_variable_116_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_116 = value_check_109_to_variable[17:12];
assign enable_check_109_to_variable_116 = enable_check_109_to_variable[2];
// 对变量节点116传递过来的值进行组合
assign value_variable_to_check_109[17:12] = value_variable_116_to_check_109;
assign enable_variable_to_check_109[2] = enable_variable_116_to_check_109;

// 拆分后校验节点109传递给变量节点154的值以及对变量节点154传递过来的值
wire [5:0] value_check_109_to_variable_154;
wire enable_check_109_to_variable_154;
wire [5:0] value_variable_154_to_check_109;
wire enable_variable_154_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_154 = value_check_109_to_variable[23:18];
assign enable_check_109_to_variable_154 = enable_check_109_to_variable[3];
// 对变量节点154传递过来的值进行组合
assign value_variable_to_check_109[23:18] = value_variable_154_to_check_109;
assign enable_variable_to_check_109[3] = enable_variable_154_to_check_109;

// 拆分后校验节点109传递给变量节点184的值以及对变量节点184传递过来的值
wire [5:0] value_check_109_to_variable_184;
wire enable_check_109_to_variable_184;
wire [5:0] value_variable_184_to_check_109;
wire enable_variable_184_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_184 = value_check_109_to_variable[29:24];
assign enable_check_109_to_variable_184 = enable_check_109_to_variable[4];
// 对变量节点184传递过来的值进行组合
assign value_variable_to_check_109[29:24] = value_variable_184_to_check_109;
assign enable_variable_to_check_109[4] = enable_variable_184_to_check_109;

// 拆分后校验节点109传递给变量节点236的值以及对变量节点236传递过来的值
wire [5:0] value_check_109_to_variable_236;
wire enable_check_109_to_variable_236;
wire [5:0] value_variable_236_to_check_109;
wire enable_variable_236_to_check_109;
// 对校验节点109的输出值进行拆分
assign value_check_109_to_variable_236 = value_check_109_to_variable[35:30];
assign enable_check_109_to_variable_236 = enable_check_109_to_variable[5];
// 对变量节点236传递过来的值进行组合
assign value_variable_to_check_109[35:30] = value_variable_236_to_check_109;
assign enable_variable_to_check_109[5] = enable_variable_236_to_check_109;


// 校验节点110的接口
wire [35:0] value_variable_to_check_110;
wire [35:0] value_check_110_to_variable;
wire [5:0] enable_variable_to_check_110;
wire [5:0] enable_check_110_to_variable;

// 拆分后校验节点110传递给变量节点27的值以及对变量节点27传递过来的值
wire [5:0] value_check_110_to_variable_27;
wire enable_check_110_to_variable_27;
wire [5:0] value_variable_27_to_check_110;
wire enable_variable_27_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_27 = value_check_110_to_variable[5:0];
assign enable_check_110_to_variable_27 = enable_check_110_to_variable[0];
// 对变量节点27传递过来的值进行组合
assign value_variable_to_check_110[5:0] = value_variable_27_to_check_110;
assign enable_variable_to_check_110[0] = enable_variable_27_to_check_110;

// 拆分后校验节点110传递给变量节点53的值以及对变量节点53传递过来的值
wire [5:0] value_check_110_to_variable_53;
wire enable_check_110_to_variable_53;
wire [5:0] value_variable_53_to_check_110;
wire enable_variable_53_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_53 = value_check_110_to_variable[11:6];
assign enable_check_110_to_variable_53 = enable_check_110_to_variable[1];
// 对变量节点53传递过来的值进行组合
assign value_variable_to_check_110[11:6] = value_variable_53_to_check_110;
assign enable_variable_to_check_110[1] = enable_variable_53_to_check_110;

// 拆分后校验节点110传递给变量节点84的值以及对变量节点84传递过来的值
wire [5:0] value_check_110_to_variable_84;
wire enable_check_110_to_variable_84;
wire [5:0] value_variable_84_to_check_110;
wire enable_variable_84_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_84 = value_check_110_to_variable[17:12];
assign enable_check_110_to_variable_84 = enable_check_110_to_variable[2];
// 对变量节点84传递过来的值进行组合
assign value_variable_to_check_110[17:12] = value_variable_84_to_check_110;
assign enable_variable_to_check_110[2] = enable_variable_84_to_check_110;

// 拆分后校验节点110传递给变量节点171的值以及对变量节点171传递过来的值
wire [5:0] value_check_110_to_variable_171;
wire enable_check_110_to_variable_171;
wire [5:0] value_variable_171_to_check_110;
wire enable_variable_171_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_171 = value_check_110_to_variable[23:18];
assign enable_check_110_to_variable_171 = enable_check_110_to_variable[3];
// 对变量节点171传递过来的值进行组合
assign value_variable_to_check_110[23:18] = value_variable_171_to_check_110;
assign enable_variable_to_check_110[3] = enable_variable_171_to_check_110;

// 拆分后校验节点110传递给变量节点206的值以及对变量节点206传递过来的值
wire [5:0] value_check_110_to_variable_206;
wire enable_check_110_to_variable_206;
wire [5:0] value_variable_206_to_check_110;
wire enable_variable_206_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_206 = value_check_110_to_variable[29:24];
assign enable_check_110_to_variable_206 = enable_check_110_to_variable[4];
// 对变量节点206传递过来的值进行组合
assign value_variable_to_check_110[29:24] = value_variable_206_to_check_110;
assign enable_variable_to_check_110[4] = enable_variable_206_to_check_110;

// 拆分后校验节点110传递给变量节点241的值以及对变量节点241传递过来的值
wire [5:0] value_check_110_to_variable_241;
wire enable_check_110_to_variable_241;
wire [5:0] value_variable_241_to_check_110;
wire enable_variable_241_to_check_110;
// 对校验节点110的输出值进行拆分
assign value_check_110_to_variable_241 = value_check_110_to_variable[35:30];
assign enable_check_110_to_variable_241 = enable_check_110_to_variable[5];
// 对变量节点241传递过来的值进行组合
assign value_variable_to_check_110[35:30] = value_variable_241_to_check_110;
assign enable_variable_to_check_110[5] = enable_variable_241_to_check_110;


// 校验节点111的接口
wire [35:0] value_variable_to_check_111;
wire [35:0] value_check_111_to_variable;
wire [5:0] enable_variable_to_check_111;
wire [5:0] enable_check_111_to_variable;

// 拆分后校验节点111传递给变量节点10的值以及对变量节点10传递过来的值
wire [5:0] value_check_111_to_variable_10;
wire enable_check_111_to_variable_10;
wire [5:0] value_variable_10_to_check_111;
wire enable_variable_10_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_10 = value_check_111_to_variable[5:0];
assign enable_check_111_to_variable_10 = enable_check_111_to_variable[0];
// 对变量节点10传递过来的值进行组合
assign value_variable_to_check_111[5:0] = value_variable_10_to_check_111;
assign enable_variable_to_check_111[0] = enable_variable_10_to_check_111;

// 拆分后校验节点111传递给变量节点74的值以及对变量节点74传递过来的值
wire [5:0] value_check_111_to_variable_74;
wire enable_check_111_to_variable_74;
wire [5:0] value_variable_74_to_check_111;
wire enable_variable_74_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_74 = value_check_111_to_variable[11:6];
assign enable_check_111_to_variable_74 = enable_check_111_to_variable[1];
// 对变量节点74传递过来的值进行组合
assign value_variable_to_check_111[11:6] = value_variable_74_to_check_111;
assign enable_variable_to_check_111[1] = enable_variable_74_to_check_111;

// 拆分后校验节点111传递给变量节点108的值以及对变量节点108传递过来的值
wire [5:0] value_check_111_to_variable_108;
wire enable_check_111_to_variable_108;
wire [5:0] value_variable_108_to_check_111;
wire enable_variable_108_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_108 = value_check_111_to_variable[17:12];
assign enable_check_111_to_variable_108 = enable_check_111_to_variable[2];
// 对变量节点108传递过来的值进行组合
assign value_variable_to_check_111[17:12] = value_variable_108_to_check_111;
assign enable_variable_to_check_111[2] = enable_variable_108_to_check_111;

// 拆分后校验节点111传递给变量节点153的值以及对变量节点153传递过来的值
wire [5:0] value_check_111_to_variable_153;
wire enable_check_111_to_variable_153;
wire [5:0] value_variable_153_to_check_111;
wire enable_variable_153_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_153 = value_check_111_to_variable[23:18];
assign enable_check_111_to_variable_153 = enable_check_111_to_variable[3];
// 对变量节点153传递过来的值进行组合
assign value_variable_to_check_111[23:18] = value_variable_153_to_check_111;
assign enable_variable_to_check_111[3] = enable_variable_153_to_check_111;

// 拆分后校验节点111传递给变量节点187的值以及对变量节点187传递过来的值
wire [5:0] value_check_111_to_variable_187;
wire enable_check_111_to_variable_187;
wire [5:0] value_variable_187_to_check_111;
wire enable_variable_187_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_187 = value_check_111_to_variable[29:24];
assign enable_check_111_to_variable_187 = enable_check_111_to_variable[4];
// 对变量节点187传递过来的值进行组合
assign value_variable_to_check_111[29:24] = value_variable_187_to_check_111;
assign enable_variable_to_check_111[4] = enable_variable_187_to_check_111;

// 拆分后校验节点111传递给变量节点255的值以及对变量节点255传递过来的值
wire [5:0] value_check_111_to_variable_255;
wire enable_check_111_to_variable_255;
wire [5:0] value_variable_255_to_check_111;
wire enable_variable_255_to_check_111;
// 对校验节点111的输出值进行拆分
assign value_check_111_to_variable_255 = value_check_111_to_variable[35:30];
assign enable_check_111_to_variable_255 = enable_check_111_to_variable[5];
// 对变量节点255传递过来的值进行组合
assign value_variable_to_check_111[35:30] = value_variable_255_to_check_111;
assign enable_variable_to_check_111[5] = enable_variable_255_to_check_111;


// 校验节点112的接口
wire [35:0] value_variable_to_check_112;
wire [35:0] value_check_112_to_variable;
wire [5:0] enable_variable_to_check_112;
wire [5:0] enable_check_112_to_variable;

// 拆分后校验节点112传递给变量节点36的值以及对变量节点36传递过来的值
wire [5:0] value_check_112_to_variable_36;
wire enable_check_112_to_variable_36;
wire [5:0] value_variable_36_to_check_112;
wire enable_variable_36_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_36 = value_check_112_to_variable[5:0];
assign enable_check_112_to_variable_36 = enable_check_112_to_variable[0];
// 对变量节点36传递过来的值进行组合
assign value_variable_to_check_112[5:0] = value_variable_36_to_check_112;
assign enable_variable_to_check_112[0] = enable_variable_36_to_check_112;

// 拆分后校验节点112传递给变量节点80的值以及对变量节点80传递过来的值
wire [5:0] value_check_112_to_variable_80;
wire enable_check_112_to_variable_80;
wire [5:0] value_variable_80_to_check_112;
wire enable_variable_80_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_80 = value_check_112_to_variable[11:6];
assign enable_check_112_to_variable_80 = enable_check_112_to_variable[1];
// 对变量节点80传递过来的值进行组合
assign value_variable_to_check_112[11:6] = value_variable_80_to_check_112;
assign enable_variable_to_check_112[1] = enable_variable_80_to_check_112;

// 拆分后校验节点112传递给变量节点91的值以及对变量节点91传递过来的值
wire [5:0] value_check_112_to_variable_91;
wire enable_check_112_to_variable_91;
wire [5:0] value_variable_91_to_check_112;
wire enable_variable_91_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_91 = value_check_112_to_variable[17:12];
assign enable_check_112_to_variable_91 = enable_check_112_to_variable[2];
// 对变量节点91传递过来的值进行组合
assign value_variable_to_check_112[17:12] = value_variable_91_to_check_112;
assign enable_variable_to_check_112[2] = enable_variable_91_to_check_112;

// 拆分后校验节点112传递给变量节点145的值以及对变量节点145传递过来的值
wire [5:0] value_check_112_to_variable_145;
wire enable_check_112_to_variable_145;
wire [5:0] value_variable_145_to_check_112;
wire enable_variable_145_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_145 = value_check_112_to_variable[23:18];
assign enable_check_112_to_variable_145 = enable_check_112_to_variable[3];
// 对变量节点145传递过来的值进行组合
assign value_variable_to_check_112[23:18] = value_variable_145_to_check_112;
assign enable_variable_to_check_112[3] = enable_variable_145_to_check_112;

// 拆分后校验节点112传递给变量节点178的值以及对变量节点178传递过来的值
wire [5:0] value_check_112_to_variable_178;
wire enable_check_112_to_variable_178;
wire [5:0] value_variable_178_to_check_112;
wire enable_variable_178_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_178 = value_check_112_to_variable[29:24];
assign enable_check_112_to_variable_178 = enable_check_112_to_variable[4];
// 对变量节点178传递过来的值进行组合
assign value_variable_to_check_112[29:24] = value_variable_178_to_check_112;
assign enable_variable_to_check_112[4] = enable_variable_178_to_check_112;

// 拆分后校验节点112传递给变量节点241的值以及对变量节点241传递过来的值
wire [5:0] value_check_112_to_variable_241;
wire enable_check_112_to_variable_241;
wire [5:0] value_variable_241_to_check_112;
wire enable_variable_241_to_check_112;
// 对校验节点112的输出值进行拆分
assign value_check_112_to_variable_241 = value_check_112_to_variable[35:30];
assign enable_check_112_to_variable_241 = enable_check_112_to_variable[5];
// 对变量节点241传递过来的值进行组合
assign value_variable_to_check_112[35:30] = value_variable_241_to_check_112;
assign enable_variable_to_check_112[5] = enable_variable_241_to_check_112;


// 校验节点113的接口
wire [35:0] value_variable_to_check_113;
wire [35:0] value_check_113_to_variable;
wire [5:0] enable_variable_to_check_113;
wire [5:0] enable_check_113_to_variable;

// 拆分后校验节点113传递给变量节点26的值以及对变量节点26传递过来的值
wire [5:0] value_check_113_to_variable_26;
wire enable_check_113_to_variable_26;
wire [5:0] value_variable_26_to_check_113;
wire enable_variable_26_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_26 = value_check_113_to_variable[5:0];
assign enable_check_113_to_variable_26 = enable_check_113_to_variable[0];
// 对变量节点26传递过来的值进行组合
assign value_variable_to_check_113[5:0] = value_variable_26_to_check_113;
assign enable_variable_to_check_113[0] = enable_variable_26_to_check_113;

// 拆分后校验节点113传递给变量节点69的值以及对变量节点69传递过来的值
wire [5:0] value_check_113_to_variable_69;
wire enable_check_113_to_variable_69;
wire [5:0] value_variable_69_to_check_113;
wire enable_variable_69_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_69 = value_check_113_to_variable[11:6];
assign enable_check_113_to_variable_69 = enable_check_113_to_variable[1];
// 对变量节点69传递过来的值进行组合
assign value_variable_to_check_113[11:6] = value_variable_69_to_check_113;
assign enable_variable_to_check_113[1] = enable_variable_69_to_check_113;

// 拆分后校验节点113传递给变量节点107的值以及对变量节点107传递过来的值
wire [5:0] value_check_113_to_variable_107;
wire enable_check_113_to_variable_107;
wire [5:0] value_variable_107_to_check_113;
wire enable_variable_107_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_107 = value_check_113_to_variable[17:12];
assign enable_check_113_to_variable_107 = enable_check_113_to_variable[2];
// 对变量节点107传递过来的值进行组合
assign value_variable_to_check_113[17:12] = value_variable_107_to_check_113;
assign enable_variable_to_check_113[2] = enable_variable_107_to_check_113;

// 拆分后校验节点113传递给变量节点163的值以及对变量节点163传递过来的值
wire [5:0] value_check_113_to_variable_163;
wire enable_check_113_to_variable_163;
wire [5:0] value_variable_163_to_check_113;
wire enable_variable_163_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_163 = value_check_113_to_variable[23:18];
assign enable_check_113_to_variable_163 = enable_check_113_to_variable[3];
// 对变量节点163传递过来的值进行组合
assign value_variable_to_check_113[23:18] = value_variable_163_to_check_113;
assign enable_variable_to_check_113[3] = enable_variable_163_to_check_113;

// 拆分后校验节点113传递给变量节点213的值以及对变量节点213传递过来的值
wire [5:0] value_check_113_to_variable_213;
wire enable_check_113_to_variable_213;
wire [5:0] value_variable_213_to_check_113;
wire enable_variable_213_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_213 = value_check_113_to_variable[29:24];
assign enable_check_113_to_variable_213 = enable_check_113_to_variable[4];
// 对变量节点213传递过来的值进行组合
assign value_variable_to_check_113[29:24] = value_variable_213_to_check_113;
assign enable_variable_to_check_113[4] = enable_variable_213_to_check_113;

// 拆分后校验节点113传递给变量节点238的值以及对变量节点238传递过来的值
wire [5:0] value_check_113_to_variable_238;
wire enable_check_113_to_variable_238;
wire [5:0] value_variable_238_to_check_113;
wire enable_variable_238_to_check_113;
// 对校验节点113的输出值进行拆分
assign value_check_113_to_variable_238 = value_check_113_to_variable[35:30];
assign enable_check_113_to_variable_238 = enable_check_113_to_variable[5];
// 对变量节点238传递过来的值进行组合
assign value_variable_to_check_113[35:30] = value_variable_238_to_check_113;
assign enable_variable_to_check_113[5] = enable_variable_238_to_check_113;


// 校验节点114的接口
wire [35:0] value_variable_to_check_114;
wire [35:0] value_check_114_to_variable;
wire [5:0] enable_variable_to_check_114;
wire [5:0] enable_check_114_to_variable;

// 拆分后校验节点114传递给变量节点5的值以及对变量节点5传递过来的值
wire [5:0] value_check_114_to_variable_5;
wire enable_check_114_to_variable_5;
wire [5:0] value_variable_5_to_check_114;
wire enable_variable_5_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_5 = value_check_114_to_variable[5:0];
assign enable_check_114_to_variable_5 = enable_check_114_to_variable[0];
// 对变量节点5传递过来的值进行组合
assign value_variable_to_check_114[5:0] = value_variable_5_to_check_114;
assign enable_variable_to_check_114[0] = enable_variable_5_to_check_114;

// 拆分后校验节点114传递给变量节点85的值以及对变量节点85传递过来的值
wire [5:0] value_check_114_to_variable_85;
wire enable_check_114_to_variable_85;
wire [5:0] value_variable_85_to_check_114;
wire enable_variable_85_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_85 = value_check_114_to_variable[11:6];
assign enable_check_114_to_variable_85 = enable_check_114_to_variable[1];
// 对变量节点85传递过来的值进行组合
assign value_variable_to_check_114[11:6] = value_variable_85_to_check_114;
assign enable_variable_to_check_114[1] = enable_variable_85_to_check_114;

// 拆分后校验节点114传递给变量节点120的值以及对变量节点120传递过来的值
wire [5:0] value_check_114_to_variable_120;
wire enable_check_114_to_variable_120;
wire [5:0] value_variable_120_to_check_114;
wire enable_variable_120_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_120 = value_check_114_to_variable[17:12];
assign enable_check_114_to_variable_120 = enable_check_114_to_variable[2];
// 对变量节点120传递过来的值进行组合
assign value_variable_to_check_114[17:12] = value_variable_120_to_check_114;
assign enable_variable_to_check_114[2] = enable_variable_120_to_check_114;

// 拆分后校验节点114传递给变量节点168的值以及对变量节点168传递过来的值
wire [5:0] value_check_114_to_variable_168;
wire enable_check_114_to_variable_168;
wire [5:0] value_variable_168_to_check_114;
wire enable_variable_168_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_168 = value_check_114_to_variable[23:18];
assign enable_check_114_to_variable_168 = enable_check_114_to_variable[3];
// 对变量节点168传递过来的值进行组合
assign value_variable_to_check_114[23:18] = value_variable_168_to_check_114;
assign enable_variable_to_check_114[3] = enable_variable_168_to_check_114;

// 拆分后校验节点114传递给变量节点211的值以及对变量节点211传递过来的值
wire [5:0] value_check_114_to_variable_211;
wire enable_check_114_to_variable_211;
wire [5:0] value_variable_211_to_check_114;
wire enable_variable_211_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_211 = value_check_114_to_variable[29:24];
assign enable_check_114_to_variable_211 = enable_check_114_to_variable[4];
// 对变量节点211传递过来的值进行组合
assign value_variable_to_check_114[29:24] = value_variable_211_to_check_114;
assign enable_variable_to_check_114[4] = enable_variable_211_to_check_114;

// 拆分后校验节点114传递给变量节点253的值以及对变量节点253传递过来的值
wire [5:0] value_check_114_to_variable_253;
wire enable_check_114_to_variable_253;
wire [5:0] value_variable_253_to_check_114;
wire enable_variable_253_to_check_114;
// 对校验节点114的输出值进行拆分
assign value_check_114_to_variable_253 = value_check_114_to_variable[35:30];
assign enable_check_114_to_variable_253 = enable_check_114_to_variable[5];
// 对变量节点253传递过来的值进行组合
assign value_variable_to_check_114[35:30] = value_variable_253_to_check_114;
assign enable_variable_to_check_114[5] = enable_variable_253_to_check_114;


// 校验节点115的接口
wire [35:0] value_variable_to_check_115;
wire [35:0] value_check_115_to_variable;
wire [5:0] enable_variable_to_check_115;
wire [5:0] enable_check_115_to_variable;

// 拆分后校验节点115传递给变量节点42的值以及对变量节点42传递过来的值
wire [5:0] value_check_115_to_variable_42;
wire enable_check_115_to_variable_42;
wire [5:0] value_variable_42_to_check_115;
wire enable_variable_42_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_42 = value_check_115_to_variable[5:0];
assign enable_check_115_to_variable_42 = enable_check_115_to_variable[0];
// 对变量节点42传递过来的值进行组合
assign value_variable_to_check_115[5:0] = value_variable_42_to_check_115;
assign enable_variable_to_check_115[0] = enable_variable_42_to_check_115;

// 拆分后校验节点115传递给变量节点69的值以及对变量节点69传递过来的值
wire [5:0] value_check_115_to_variable_69;
wire enable_check_115_to_variable_69;
wire [5:0] value_variable_69_to_check_115;
wire enable_variable_69_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_69 = value_check_115_to_variable[11:6];
assign enable_check_115_to_variable_69 = enable_check_115_to_variable[1];
// 对变量节点69传递过来的值进行组合
assign value_variable_to_check_115[11:6] = value_variable_69_to_check_115;
assign enable_variable_to_check_115[1] = enable_variable_69_to_check_115;

// 拆分后校验节点115传递给变量节点123的值以及对变量节点123传递过来的值
wire [5:0] value_check_115_to_variable_123;
wire enable_check_115_to_variable_123;
wire [5:0] value_variable_123_to_check_115;
wire enable_variable_123_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_123 = value_check_115_to_variable[17:12];
assign enable_check_115_to_variable_123 = enable_check_115_to_variable[2];
// 对变量节点123传递过来的值进行组合
assign value_variable_to_check_115[17:12] = value_variable_123_to_check_115;
assign enable_variable_to_check_115[2] = enable_variable_123_to_check_115;

// 拆分后校验节点115传递给变量节点159的值以及对变量节点159传递过来的值
wire [5:0] value_check_115_to_variable_159;
wire enable_check_115_to_variable_159;
wire [5:0] value_variable_159_to_check_115;
wire enable_variable_159_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_159 = value_check_115_to_variable[23:18];
assign enable_check_115_to_variable_159 = enable_check_115_to_variable[3];
// 对变量节点159传递过来的值进行组合
assign value_variable_to_check_115[23:18] = value_variable_159_to_check_115;
assign enable_variable_to_check_115[3] = enable_variable_159_to_check_115;

// 拆分后校验节点115传递给变量节点194的值以及对变量节点194传递过来的值
wire [5:0] value_check_115_to_variable_194;
wire enable_check_115_to_variable_194;
wire [5:0] value_variable_194_to_check_115;
wire enable_variable_194_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_194 = value_check_115_to_variable[29:24];
assign enable_check_115_to_variable_194 = enable_check_115_to_variable[4];
// 对变量节点194传递过来的值进行组合
assign value_variable_to_check_115[29:24] = value_variable_194_to_check_115;
assign enable_variable_to_check_115[4] = enable_variable_194_to_check_115;

// 拆分后校验节点115传递给变量节点251的值以及对变量节点251传递过来的值
wire [5:0] value_check_115_to_variable_251;
wire enable_check_115_to_variable_251;
wire [5:0] value_variable_251_to_check_115;
wire enable_variable_251_to_check_115;
// 对校验节点115的输出值进行拆分
assign value_check_115_to_variable_251 = value_check_115_to_variable[35:30];
assign enable_check_115_to_variable_251 = enable_check_115_to_variable[5];
// 对变量节点251传递过来的值进行组合
assign value_variable_to_check_115[35:30] = value_variable_251_to_check_115;
assign enable_variable_to_check_115[5] = enable_variable_251_to_check_115;


// 校验节点116的接口
wire [35:0] value_variable_to_check_116;
wire [35:0] value_check_116_to_variable;
wire [5:0] enable_variable_to_check_116;
wire [5:0] enable_check_116_to_variable;

// 拆分后校验节点116传递给变量节点25的值以及对变量节点25传递过来的值
wire [5:0] value_check_116_to_variable_25;
wire enable_check_116_to_variable_25;
wire [5:0] value_variable_25_to_check_116;
wire enable_variable_25_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_25 = value_check_116_to_variable[5:0];
assign enable_check_116_to_variable_25 = enable_check_116_to_variable[0];
// 对变量节点25传递过来的值进行组合
assign value_variable_to_check_116[5:0] = value_variable_25_to_check_116;
assign enable_variable_to_check_116[0] = enable_variable_25_to_check_116;

// 拆分后校验节点116传递给变量节点66的值以及对变量节点66传递过来的值
wire [5:0] value_check_116_to_variable_66;
wire enable_check_116_to_variable_66;
wire [5:0] value_variable_66_to_check_116;
wire enable_variable_66_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_66 = value_check_116_to_variable[11:6];
assign enable_check_116_to_variable_66 = enable_check_116_to_variable[1];
// 对变量节点66传递过来的值进行组合
assign value_variable_to_check_116[11:6] = value_variable_66_to_check_116;
assign enable_variable_to_check_116[1] = enable_variable_66_to_check_116;

// 拆分后校验节点116传递给变量节点121的值以及对变量节点121传递过来的值
wire [5:0] value_check_116_to_variable_121;
wire enable_check_116_to_variable_121;
wire [5:0] value_variable_121_to_check_116;
wire enable_variable_121_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_121 = value_check_116_to_variable[17:12];
assign enable_check_116_to_variable_121 = enable_check_116_to_variable[2];
// 对变量节点121传递过来的值进行组合
assign value_variable_to_check_116[17:12] = value_variable_121_to_check_116;
assign enable_variable_to_check_116[2] = enable_variable_121_to_check_116;

// 拆分后校验节点116传递给变量节点170的值以及对变量节点170传递过来的值
wire [5:0] value_check_116_to_variable_170;
wire enable_check_116_to_variable_170;
wire [5:0] value_variable_170_to_check_116;
wire enable_variable_170_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_170 = value_check_116_to_variable[23:18];
assign enable_check_116_to_variable_170 = enable_check_116_to_variable[3];
// 对变量节点170传递过来的值进行组合
assign value_variable_to_check_116[23:18] = value_variable_170_to_check_116;
assign enable_variable_to_check_116[3] = enable_variable_170_to_check_116;

// 拆分后校验节点116传递给变量节点198的值以及对变量节点198传递过来的值
wire [5:0] value_check_116_to_variable_198;
wire enable_check_116_to_variable_198;
wire [5:0] value_variable_198_to_check_116;
wire enable_variable_198_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_198 = value_check_116_to_variable[29:24];
assign enable_check_116_to_variable_198 = enable_check_116_to_variable[4];
// 对变量节点198传递过来的值进行组合
assign value_variable_to_check_116[29:24] = value_variable_198_to_check_116;
assign enable_variable_to_check_116[4] = enable_variable_198_to_check_116;

// 拆分后校验节点116传递给变量节点224的值以及对变量节点224传递过来的值
wire [5:0] value_check_116_to_variable_224;
wire enable_check_116_to_variable_224;
wire [5:0] value_variable_224_to_check_116;
wire enable_variable_224_to_check_116;
// 对校验节点116的输出值进行拆分
assign value_check_116_to_variable_224 = value_check_116_to_variable[35:30];
assign enable_check_116_to_variable_224 = enable_check_116_to_variable[5];
// 对变量节点224传递过来的值进行组合
assign value_variable_to_check_116[35:30] = value_variable_224_to_check_116;
assign enable_variable_to_check_116[5] = enable_variable_224_to_check_116;


// 校验节点117的接口
wire [35:0] value_variable_to_check_117;
wire [35:0] value_check_117_to_variable;
wire [5:0] enable_variable_to_check_117;
wire [5:0] enable_check_117_to_variable;

// 拆分后校验节点117传递给变量节点11的值以及对变量节点11传递过来的值
wire [5:0] value_check_117_to_variable_11;
wire enable_check_117_to_variable_11;
wire [5:0] value_variable_11_to_check_117;
wire enable_variable_11_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_11 = value_check_117_to_variable[5:0];
assign enable_check_117_to_variable_11 = enable_check_117_to_variable[0];
// 对变量节点11传递过来的值进行组合
assign value_variable_to_check_117[5:0] = value_variable_11_to_check_117;
assign enable_variable_to_check_117[0] = enable_variable_11_to_check_117;

// 拆分后校验节点117传递给变量节点56的值以及对变量节点56传递过来的值
wire [5:0] value_check_117_to_variable_56;
wire enable_check_117_to_variable_56;
wire [5:0] value_variable_56_to_check_117;
wire enable_variable_56_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_56 = value_check_117_to_variable[11:6];
assign enable_check_117_to_variable_56 = enable_check_117_to_variable[1];
// 对变量节点56传递过来的值进行组合
assign value_variable_to_check_117[11:6] = value_variable_56_to_check_117;
assign enable_variable_to_check_117[1] = enable_variable_56_to_check_117;

// 拆分后校验节点117传递给变量节点130的值以及对变量节点130传递过来的值
wire [5:0] value_check_117_to_variable_130;
wire enable_check_117_to_variable_130;
wire [5:0] value_variable_130_to_check_117;
wire enable_variable_130_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_130 = value_check_117_to_variable[17:12];
assign enable_check_117_to_variable_130 = enable_check_117_to_variable[2];
// 对变量节点130传递过来的值进行组合
assign value_variable_to_check_117[17:12] = value_variable_130_to_check_117;
assign enable_variable_to_check_117[2] = enable_variable_130_to_check_117;

// 拆分后校验节点117传递给变量节点142的值以及对变量节点142传递过来的值
wire [5:0] value_check_117_to_variable_142;
wire enable_check_117_to_variable_142;
wire [5:0] value_variable_142_to_check_117;
wire enable_variable_142_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_142 = value_check_117_to_variable[23:18];
assign enable_check_117_to_variable_142 = enable_check_117_to_variable[3];
// 对变量节点142传递过来的值进行组合
assign value_variable_to_check_117[23:18] = value_variable_142_to_check_117;
assign enable_variable_to_check_117[3] = enable_variable_142_to_check_117;

// 拆分后校验节点117传递给变量节点179的值以及对变量节点179传递过来的值
wire [5:0] value_check_117_to_variable_179;
wire enable_check_117_to_variable_179;
wire [5:0] value_variable_179_to_check_117;
wire enable_variable_179_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_179 = value_check_117_to_variable[29:24];
assign enable_check_117_to_variable_179 = enable_check_117_to_variable[4];
// 对变量节点179传递过来的值进行组合
assign value_variable_to_check_117[29:24] = value_variable_179_to_check_117;
assign enable_variable_to_check_117[4] = enable_variable_179_to_check_117;

// 拆分后校验节点117传递给变量节点214的值以及对变量节点214传递过来的值
wire [5:0] value_check_117_to_variable_214;
wire enable_check_117_to_variable_214;
wire [5:0] value_variable_214_to_check_117;
wire enable_variable_214_to_check_117;
// 对校验节点117的输出值进行拆分
assign value_check_117_to_variable_214 = value_check_117_to_variable[35:30];
assign enable_check_117_to_variable_214 = enable_check_117_to_variable[5];
// 对变量节点214传递过来的值进行组合
assign value_variable_to_check_117[35:30] = value_variable_214_to_check_117;
assign enable_variable_to_check_117[5] = enable_variable_214_to_check_117;


// 校验节点118的接口
wire [35:0] value_variable_to_check_118;
wire [35:0] value_check_118_to_variable;
wire [5:0] enable_variable_to_check_118;
wire [5:0] enable_check_118_to_variable;

// 拆分后校验节点118传递给变量节点39的值以及对变量节点39传递过来的值
wire [5:0] value_check_118_to_variable_39;
wire enable_check_118_to_variable_39;
wire [5:0] value_variable_39_to_check_118;
wire enable_variable_39_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_39 = value_check_118_to_variable[5:0];
assign enable_check_118_to_variable_39 = enable_check_118_to_variable[0];
// 对变量节点39传递过来的值进行组合
assign value_variable_to_check_118[5:0] = value_variable_39_to_check_118;
assign enable_variable_to_check_118[0] = enable_variable_39_to_check_118;

// 拆分后校验节点118传递给变量节点70的值以及对变量节点70传递过来的值
wire [5:0] value_check_118_to_variable_70;
wire enable_check_118_to_variable_70;
wire [5:0] value_variable_70_to_check_118;
wire enable_variable_70_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_70 = value_check_118_to_variable[11:6];
assign enable_check_118_to_variable_70 = enable_check_118_to_variable[1];
// 对变量节点70传递过来的值进行组合
assign value_variable_to_check_118[11:6] = value_variable_70_to_check_118;
assign enable_variable_to_check_118[1] = enable_variable_70_to_check_118;

// 拆分后校验节点118传递给变量节点93的值以及对变量节点93传递过来的值
wire [5:0] value_check_118_to_variable_93;
wire enable_check_118_to_variable_93;
wire [5:0] value_variable_93_to_check_118;
wire enable_variable_93_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_93 = value_check_118_to_variable[17:12];
assign enable_check_118_to_variable_93 = enable_check_118_to_variable[2];
// 对变量节点93传递过来的值进行组合
assign value_variable_to_check_118[17:12] = value_variable_93_to_check_118;
assign enable_variable_to_check_118[2] = enable_variable_93_to_check_118;

// 拆分后校验节点118传递给变量节点134的值以及对变量节点134传递过来的值
wire [5:0] value_check_118_to_variable_134;
wire enable_check_118_to_variable_134;
wire [5:0] value_variable_134_to_check_118;
wire enable_variable_134_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_134 = value_check_118_to_variable[23:18];
assign enable_check_118_to_variable_134 = enable_check_118_to_variable[3];
// 对变量节点134传递过来的值进行组合
assign value_variable_to_check_118[23:18] = value_variable_134_to_check_118;
assign enable_variable_to_check_118[3] = enable_variable_134_to_check_118;

// 拆分后校验节点118传递给变量节点152的值以及对变量节点152传递过来的值
wire [5:0] value_check_118_to_variable_152;
wire enable_check_118_to_variable_152;
wire [5:0] value_variable_152_to_check_118;
wire enable_variable_152_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_152 = value_check_118_to_variable[29:24];
assign enable_check_118_to_variable_152 = enable_check_118_to_variable[4];
// 对变量节点152传递过来的值进行组合
assign value_variable_to_check_118[29:24] = value_variable_152_to_check_118;
assign enable_variable_to_check_118[4] = enable_variable_152_to_check_118;

// 拆分后校验节点118传递给变量节点252的值以及对变量节点252传递过来的值
wire [5:0] value_check_118_to_variable_252;
wire enable_check_118_to_variable_252;
wire [5:0] value_variable_252_to_check_118;
wire enable_variable_252_to_check_118;
// 对校验节点118的输出值进行拆分
assign value_check_118_to_variable_252 = value_check_118_to_variable[35:30];
assign enable_check_118_to_variable_252 = enable_check_118_to_variable[5];
// 对变量节点252传递过来的值进行组合
assign value_variable_to_check_118[35:30] = value_variable_252_to_check_118;
assign enable_variable_to_check_118[5] = enable_variable_252_to_check_118;


// 校验节点119的接口
wire [35:0] value_variable_to_check_119;
wire [35:0] value_check_119_to_variable;
wire [5:0] enable_variable_to_check_119;
wire [5:0] enable_check_119_to_variable;

// 拆分后校验节点119传递给变量节点12的值以及对变量节点12传递过来的值
wire [5:0] value_check_119_to_variable_12;
wire enable_check_119_to_variable_12;
wire [5:0] value_variable_12_to_check_119;
wire enable_variable_12_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_12 = value_check_119_to_variable[5:0];
assign enable_check_119_to_variable_12 = enable_check_119_to_variable[0];
// 对变量节点12传递过来的值进行组合
assign value_variable_to_check_119[5:0] = value_variable_12_to_check_119;
assign enable_variable_to_check_119[0] = enable_variable_12_to_check_119;

// 拆分后校验节点119传递给变量节点79的值以及对变量节点79传递过来的值
wire [5:0] value_check_119_to_variable_79;
wire enable_check_119_to_variable_79;
wire [5:0] value_variable_79_to_check_119;
wire enable_variable_79_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_79 = value_check_119_to_variable[11:6];
assign enable_check_119_to_variable_79 = enable_check_119_to_variable[1];
// 对变量节点79传递过来的值进行组合
assign value_variable_to_check_119[11:6] = value_variable_79_to_check_119;
assign enable_variable_to_check_119[1] = enable_variable_79_to_check_119;

// 拆分后校验节点119传递给变量节点105的值以及对变量节点105传递过来的值
wire [5:0] value_check_119_to_variable_105;
wire enable_check_119_to_variable_105;
wire [5:0] value_variable_105_to_check_119;
wire enable_variable_105_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_105 = value_check_119_to_variable[17:12];
assign enable_check_119_to_variable_105 = enable_check_119_to_variable[2];
// 对变量节点105传递过来的值进行组合
assign value_variable_to_check_119[17:12] = value_variable_105_to_check_119;
assign enable_variable_to_check_119[2] = enable_variable_105_to_check_119;

// 拆分后校验节点119传递给变量节点172的值以及对变量节点172传递过来的值
wire [5:0] value_check_119_to_variable_172;
wire enable_check_119_to_variable_172;
wire [5:0] value_variable_172_to_check_119;
wire enable_variable_172_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_172 = value_check_119_to_variable[23:18];
assign enable_check_119_to_variable_172 = enable_check_119_to_variable[3];
// 对变量节点172传递过来的值进行组合
assign value_variable_to_check_119[23:18] = value_variable_172_to_check_119;
assign enable_variable_to_check_119[3] = enable_variable_172_to_check_119;

// 拆分后校验节点119传递给变量节点190的值以及对变量节点190传递过来的值
wire [5:0] value_check_119_to_variable_190;
wire enable_check_119_to_variable_190;
wire [5:0] value_variable_190_to_check_119;
wire enable_variable_190_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_190 = value_check_119_to_variable[29:24];
assign enable_check_119_to_variable_190 = enable_check_119_to_variable[4];
// 对变量节点190传递过来的值进行组合
assign value_variable_to_check_119[29:24] = value_variable_190_to_check_119;
assign enable_variable_to_check_119[4] = enable_variable_190_to_check_119;

// 拆分后校验节点119传递给变量节点215的值以及对变量节点215传递过来的值
wire [5:0] value_check_119_to_variable_215;
wire enable_check_119_to_variable_215;
wire [5:0] value_variable_215_to_check_119;
wire enable_variable_215_to_check_119;
// 对校验节点119的输出值进行拆分
assign value_check_119_to_variable_215 = value_check_119_to_variable[35:30];
assign enable_check_119_to_variable_215 = enable_check_119_to_variable[5];
// 对变量节点215传递过来的值进行组合
assign value_variable_to_check_119[35:30] = value_variable_215_to_check_119;
assign enable_variable_to_check_119[5] = enable_variable_215_to_check_119;


// 校验节点120的接口
wire [35:0] value_variable_to_check_120;
wire [35:0] value_check_120_to_variable;
wire [5:0] enable_variable_to_check_120;
wire [5:0] enable_check_120_to_variable;

// 拆分后校验节点120传递给变量节点30的值以及对变量节点30传递过来的值
wire [5:0] value_check_120_to_variable_30;
wire enable_check_120_to_variable_30;
wire [5:0] value_variable_30_to_check_120;
wire enable_variable_30_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_30 = value_check_120_to_variable[5:0];
assign enable_check_120_to_variable_30 = enable_check_120_to_variable[0];
// 对变量节点30传递过来的值进行组合
assign value_variable_to_check_120[5:0] = value_variable_30_to_check_120;
assign enable_variable_to_check_120[0] = enable_variable_30_to_check_120;

// 拆分后校验节点120传递给变量节点75的值以及对变量节点75传递过来的值
wire [5:0] value_check_120_to_variable_75;
wire enable_check_120_to_variable_75;
wire [5:0] value_variable_75_to_check_120;
wire enable_variable_75_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_75 = value_check_120_to_variable[11:6];
assign enable_check_120_to_variable_75 = enable_check_120_to_variable[1];
// 对变量节点75传递过来的值进行组合
assign value_variable_to_check_120[11:6] = value_variable_75_to_check_120;
assign enable_variable_to_check_120[1] = enable_variable_75_to_check_120;

// 拆分后校验节点120传递给变量节点113的值以及对变量节点113传递过来的值
wire [5:0] value_check_120_to_variable_113;
wire enable_check_120_to_variable_113;
wire [5:0] value_variable_113_to_check_120;
wire enable_variable_113_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_113 = value_check_120_to_variable[17:12];
assign enable_check_120_to_variable_113 = enable_check_120_to_variable[2];
// 对变量节点113传递过来的值进行组合
assign value_variable_to_check_120[17:12] = value_variable_113_to_check_120;
assign enable_variable_to_check_120[2] = enable_variable_113_to_check_120;

// 拆分后校验节点120传递给变量节点157的值以及对变量节点157传递过来的值
wire [5:0] value_check_120_to_variable_157;
wire enable_check_120_to_variable_157;
wire [5:0] value_variable_157_to_check_120;
wire enable_variable_157_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_157 = value_check_120_to_variable[23:18];
assign enable_check_120_to_variable_157 = enable_check_120_to_variable[3];
// 对变量节点157传递过来的值进行组合
assign value_variable_to_check_120[23:18] = value_variable_157_to_check_120;
assign enable_variable_to_check_120[3] = enable_variable_157_to_check_120;

// 拆分后校验节点120传递给变量节点187的值以及对变量节点187传递过来的值
wire [5:0] value_check_120_to_variable_187;
wire enable_check_120_to_variable_187;
wire [5:0] value_variable_187_to_check_120;
wire enable_variable_187_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_187 = value_check_120_to_variable[29:24];
assign enable_check_120_to_variable_187 = enable_check_120_to_variable[4];
// 对变量节点187传递过来的值进行组合
assign value_variable_to_check_120[29:24] = value_variable_187_to_check_120;
assign enable_variable_to_check_120[4] = enable_variable_187_to_check_120;

// 拆分后校验节点120传递给变量节点238的值以及对变量节点238传递过来的值
wire [5:0] value_check_120_to_variable_238;
wire enable_check_120_to_variable_238;
wire [5:0] value_variable_238_to_check_120;
wire enable_variable_238_to_check_120;
// 对校验节点120的输出值进行拆分
assign value_check_120_to_variable_238 = value_check_120_to_variable[35:30];
assign enable_check_120_to_variable_238 = enable_check_120_to_variable[5];
// 对变量节点238传递过来的值进行组合
assign value_variable_to_check_120[35:30] = value_variable_238_to_check_120;
assign enable_variable_to_check_120[5] = enable_variable_238_to_check_120;


// 校验节点121的接口
wire [35:0] value_variable_to_check_121;
wire [35:0] value_check_121_to_variable;
wire [5:0] enable_variable_to_check_121;
wire [5:0] enable_check_121_to_variable;

// 拆分后校验节点121传递给变量节点16的值以及对变量节点16传递过来的值
wire [5:0] value_check_121_to_variable_16;
wire enable_check_121_to_variable_16;
wire [5:0] value_variable_16_to_check_121;
wire enable_variable_16_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_16 = value_check_121_to_variable[5:0];
assign enable_check_121_to_variable_16 = enable_check_121_to_variable[0];
// 对变量节点16传递过来的值进行组合
assign value_variable_to_check_121[5:0] = value_variable_16_to_check_121;
assign enable_variable_to_check_121[0] = enable_variable_16_to_check_121;

// 拆分后校验节点121传递给变量节点74的值以及对变量节点74传递过来的值
wire [5:0] value_check_121_to_variable_74;
wire enable_check_121_to_variable_74;
wire [5:0] value_variable_74_to_check_121;
wire enable_variable_74_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_74 = value_check_121_to_variable[11:6];
assign enable_check_121_to_variable_74 = enable_check_121_to_variable[1];
// 对变量节点74传递过来的值进行组合
assign value_variable_to_check_121[11:6] = value_variable_74_to_check_121;
assign enable_variable_to_check_121[1] = enable_variable_74_to_check_121;

// 拆分后校验节点121传递给变量节点90的值以及对变量节点90传递过来的值
wire [5:0] value_check_121_to_variable_90;
wire enable_check_121_to_variable_90;
wire [5:0] value_variable_90_to_check_121;
wire enable_variable_90_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_90 = value_check_121_to_variable[17:12];
assign enable_check_121_to_variable_90 = enable_check_121_to_variable[2];
// 对变量节点90传递过来的值进行组合
assign value_variable_to_check_121[17:12] = value_variable_90_to_check_121;
assign enable_variable_to_check_121[2] = enable_variable_90_to_check_121;

// 拆分后校验节点121传递给变量节点169的值以及对变量节点169传递过来的值
wire [5:0] value_check_121_to_variable_169;
wire enable_check_121_to_variable_169;
wire [5:0] value_variable_169_to_check_121;
wire enable_variable_169_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_169 = value_check_121_to_variable[23:18];
assign enable_check_121_to_variable_169 = enable_check_121_to_variable[3];
// 对变量节点169传递过来的值进行组合
assign value_variable_to_check_121[23:18] = value_variable_169_to_check_121;
assign enable_variable_to_check_121[3] = enable_variable_169_to_check_121;

// 拆分后校验节点121传递给变量节点209的值以及对变量节点209传递过来的值
wire [5:0] value_check_121_to_variable_209;
wire enable_check_121_to_variable_209;
wire [5:0] value_variable_209_to_check_121;
wire enable_variable_209_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_209 = value_check_121_to_variable[29:24];
assign enable_check_121_to_variable_209 = enable_check_121_to_variable[4];
// 对变量节点209传递过来的值进行组合
assign value_variable_to_check_121[29:24] = value_variable_209_to_check_121;
assign enable_variable_to_check_121[4] = enable_variable_209_to_check_121;

// 拆分后校验节点121传递给变量节点237的值以及对变量节点237传递过来的值
wire [5:0] value_check_121_to_variable_237;
wire enable_check_121_to_variable_237;
wire [5:0] value_variable_237_to_check_121;
wire enable_variable_237_to_check_121;
// 对校验节点121的输出值进行拆分
assign value_check_121_to_variable_237 = value_check_121_to_variable[35:30];
assign enable_check_121_to_variable_237 = enable_check_121_to_variable[5];
// 对变量节点237传递过来的值进行组合
assign value_variable_to_check_121[35:30] = value_variable_237_to_check_121;
assign enable_variable_to_check_121[5] = enable_variable_237_to_check_121;


// 校验节点122的接口
wire [35:0] value_variable_to_check_122;
wire [35:0] value_check_122_to_variable;
wire [5:0] enable_variable_to_check_122;
wire [5:0] enable_check_122_to_variable;

// 拆分后校验节点122传递给变量节点33的值以及对变量节点33传递过来的值
wire [5:0] value_check_122_to_variable_33;
wire enable_check_122_to_variable_33;
wire [5:0] value_variable_33_to_check_122;
wire enable_variable_33_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_33 = value_check_122_to_variable[5:0];
assign enable_check_122_to_variable_33 = enable_check_122_to_variable[0];
// 对变量节点33传递过来的值进行组合
assign value_variable_to_check_122[5:0] = value_variable_33_to_check_122;
assign enable_variable_to_check_122[0] = enable_variable_33_to_check_122;

// 拆分后校验节点122传递给变量节点51的值以及对变量节点51传递过来的值
wire [5:0] value_check_122_to_variable_51;
wire enable_check_122_to_variable_51;
wire [5:0] value_variable_51_to_check_122;
wire enable_variable_51_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_51 = value_check_122_to_variable[11:6];
assign enable_check_122_to_variable_51 = enable_check_122_to_variable[1];
// 对变量节点51传递过来的值进行组合
assign value_variable_to_check_122[11:6] = value_variable_51_to_check_122;
assign enable_variable_to_check_122[1] = enable_variable_51_to_check_122;

// 拆分后校验节点122传递给变量节点84的值以及对变量节点84传递过来的值
wire [5:0] value_check_122_to_variable_84;
wire enable_check_122_to_variable_84;
wire [5:0] value_variable_84_to_check_122;
wire enable_variable_84_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_84 = value_check_122_to_variable[17:12];
assign enable_check_122_to_variable_84 = enable_check_122_to_variable[2];
// 对变量节点84传递过来的值进行组合
assign value_variable_to_check_122[17:12] = value_variable_84_to_check_122;
assign enable_variable_to_check_122[2] = enable_variable_84_to_check_122;

// 拆分后校验节点122传递给变量节点147的值以及对变量节点147传递过来的值
wire [5:0] value_check_122_to_variable_147;
wire enable_check_122_to_variable_147;
wire [5:0] value_variable_147_to_check_122;
wire enable_variable_147_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_147 = value_check_122_to_variable[23:18];
assign enable_check_122_to_variable_147 = enable_check_122_to_variable[3];
// 对变量节点147传递过来的值进行组合
assign value_variable_to_check_122[23:18] = value_variable_147_to_check_122;
assign enable_variable_to_check_122[3] = enable_variable_147_to_check_122;

// 拆分后校验节点122传递给变量节点191的值以及对变量节点191传递过来的值
wire [5:0] value_check_122_to_variable_191;
wire enable_check_122_to_variable_191;
wire [5:0] value_variable_191_to_check_122;
wire enable_variable_191_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_191 = value_check_122_to_variable[29:24];
assign enable_check_122_to_variable_191 = enable_check_122_to_variable[4];
// 对变量节点191传递过来的值进行组合
assign value_variable_to_check_122[29:24] = value_variable_191_to_check_122;
assign enable_variable_to_check_122[4] = enable_variable_191_to_check_122;

// 拆分后校验节点122传递给变量节点255的值以及对变量节点255传递过来的值
wire [5:0] value_check_122_to_variable_255;
wire enable_check_122_to_variable_255;
wire [5:0] value_variable_255_to_check_122;
wire enable_variable_255_to_check_122;
// 对校验节点122的输出值进行拆分
assign value_check_122_to_variable_255 = value_check_122_to_variable[35:30];
assign enable_check_122_to_variable_255 = enable_check_122_to_variable[5];
// 对变量节点255传递过来的值进行组合
assign value_variable_to_check_122[35:30] = value_variable_255_to_check_122;
assign enable_variable_to_check_122[5] = enable_variable_255_to_check_122;


// 校验节点123的接口
wire [35:0] value_variable_to_check_123;
wire [35:0] value_check_123_to_variable;
wire [5:0] enable_variable_to_check_123;
wire [5:0] enable_check_123_to_variable;

// 拆分后校验节点123传递给变量节点42的值以及对变量节点42传递过来的值
wire [5:0] value_check_123_to_variable_42;
wire enable_check_123_to_variable_42;
wire [5:0] value_variable_42_to_check_123;
wire enable_variable_42_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_42 = value_check_123_to_variable[5:0];
assign enable_check_123_to_variable_42 = enable_check_123_to_variable[0];
// 对变量节点42传递过来的值进行组合
assign value_variable_to_check_123[5:0] = value_variable_42_to_check_123;
assign enable_variable_to_check_123[0] = enable_variable_42_to_check_123;

// 拆分后校验节点123传递给变量节点82的值以及对变量节点82传递过来的值
wire [5:0] value_check_123_to_variable_82;
wire enable_check_123_to_variable_82;
wire [5:0] value_variable_82_to_check_123;
wire enable_variable_82_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_82 = value_check_123_to_variable[11:6];
assign enable_check_123_to_variable_82 = enable_check_123_to_variable[1];
// 对变量节点82传递过来的值进行组合
assign value_variable_to_check_123[11:6] = value_variable_82_to_check_123;
assign enable_variable_to_check_123[1] = enable_variable_82_to_check_123;

// 拆分后校验节点123传递给变量节点100的值以及对变量节点100传递过来的值
wire [5:0] value_check_123_to_variable_100;
wire enable_check_123_to_variable_100;
wire [5:0] value_variable_100_to_check_123;
wire enable_variable_100_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_100 = value_check_123_to_variable[17:12];
assign enable_check_123_to_variable_100 = enable_check_123_to_variable[2];
// 对变量节点100传递过来的值进行组合
assign value_variable_to_check_123[17:12] = value_variable_100_to_check_123;
assign enable_variable_to_check_123[2] = enable_variable_100_to_check_123;

// 拆分后校验节点123传递给变量节点136的值以及对变量节点136传递过来的值
wire [5:0] value_check_123_to_variable_136;
wire enable_check_123_to_variable_136;
wire [5:0] value_variable_136_to_check_123;
wire enable_variable_136_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_136 = value_check_123_to_variable[23:18];
assign enable_check_123_to_variable_136 = enable_check_123_to_variable[3];
// 对变量节点136传递过来的值进行组合
assign value_variable_to_check_123[23:18] = value_variable_136_to_check_123;
assign enable_variable_to_check_123[3] = enable_variable_136_to_check_123;

// 拆分后校验节点123传递给变量节点202的值以及对变量节点202传递过来的值
wire [5:0] value_check_123_to_variable_202;
wire enable_check_123_to_variable_202;
wire [5:0] value_variable_202_to_check_123;
wire enable_variable_202_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_202 = value_check_123_to_variable[29:24];
assign enable_check_123_to_variable_202 = enable_check_123_to_variable[4];
// 对变量节点202传递过来的值进行组合
assign value_variable_to_check_123[29:24] = value_variable_202_to_check_123;
assign enable_variable_to_check_123[4] = enable_variable_202_to_check_123;

// 拆分后校验节点123传递给变量节点245的值以及对变量节点245传递过来的值
wire [5:0] value_check_123_to_variable_245;
wire enable_check_123_to_variable_245;
wire [5:0] value_variable_245_to_check_123;
wire enable_variable_245_to_check_123;
// 对校验节点123的输出值进行拆分
assign value_check_123_to_variable_245 = value_check_123_to_variable[35:30];
assign enable_check_123_to_variable_245 = enable_check_123_to_variable[5];
// 对变量节点245传递过来的值进行组合
assign value_variable_to_check_123[35:30] = value_variable_245_to_check_123;
assign enable_variable_to_check_123[5] = enable_variable_245_to_check_123;


// 校验节点124的接口
wire [35:0] value_variable_to_check_124;
wire [35:0] value_check_124_to_variable;
wire [5:0] enable_variable_to_check_124;
wire [5:0] enable_check_124_to_variable;

// 拆分后校验节点124传递给变量节点30的值以及对变量节点30传递过来的值
wire [5:0] value_check_124_to_variable_30;
wire enable_check_124_to_variable_30;
wire [5:0] value_variable_30_to_check_124;
wire enable_variable_30_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_30 = value_check_124_to_variable[5:0];
assign enable_check_124_to_variable_30 = enable_check_124_to_variable[0];
// 对变量节点30传递过来的值进行组合
assign value_variable_to_check_124[5:0] = value_variable_30_to_check_124;
assign enable_variable_to_check_124[0] = enable_variable_30_to_check_124;

// 拆分后校验节点124传递给变量节点65的值以及对变量节点65传递过来的值
wire [5:0] value_check_124_to_variable_65;
wire enable_check_124_to_variable_65;
wire [5:0] value_variable_65_to_check_124;
wire enable_variable_65_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_65 = value_check_124_to_variable[11:6];
assign enable_check_124_to_variable_65 = enable_check_124_to_variable[1];
// 对变量节点65传递过来的值进行组合
assign value_variable_to_check_124[11:6] = value_variable_65_to_check_124;
assign enable_variable_to_check_124[1] = enable_variable_65_to_check_124;

// 拆分后校验节点124传递给变量节点98的值以及对变量节点98传递过来的值
wire [5:0] value_check_124_to_variable_98;
wire enable_check_124_to_variable_98;
wire [5:0] value_variable_98_to_check_124;
wire enable_variable_98_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_98 = value_check_124_to_variable[17:12];
assign enable_check_124_to_variable_98 = enable_check_124_to_variable[2];
// 对变量节点98传递过来的值进行组合
assign value_variable_to_check_124[17:12] = value_variable_98_to_check_124;
assign enable_variable_to_check_124[2] = enable_variable_98_to_check_124;

// 拆分后校验节点124传递给变量节点167的值以及对变量节点167传递过来的值
wire [5:0] value_check_124_to_variable_167;
wire enable_check_124_to_variable_167;
wire [5:0] value_variable_167_to_check_124;
wire enable_variable_167_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_167 = value_check_124_to_variable[23:18];
assign enable_check_124_to_variable_167 = enable_check_124_to_variable[3];
// 对变量节点167传递过来的值进行组合
assign value_variable_to_check_124[23:18] = value_variable_167_to_check_124;
assign enable_variable_to_check_124[3] = enable_variable_167_to_check_124;

// 拆分后校验节点124传递给变量节点211的值以及对变量节点211传递过来的值
wire [5:0] value_check_124_to_variable_211;
wire enable_check_124_to_variable_211;
wire [5:0] value_variable_211_to_check_124;
wire enable_variable_211_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_211 = value_check_124_to_variable[29:24];
assign enable_check_124_to_variable_211 = enable_check_124_to_variable[4];
// 对变量节点211传递过来的值进行组合
assign value_variable_to_check_124[29:24] = value_variable_211_to_check_124;
assign enable_variable_to_check_124[4] = enable_variable_211_to_check_124;

// 拆分后校验节点124传递给变量节点248的值以及对变量节点248传递过来的值
wire [5:0] value_check_124_to_variable_248;
wire enable_check_124_to_variable_248;
wire [5:0] value_variable_248_to_check_124;
wire enable_variable_248_to_check_124;
// 对校验节点124的输出值进行拆分
assign value_check_124_to_variable_248 = value_check_124_to_variable[35:30];
assign enable_check_124_to_variable_248 = enable_check_124_to_variable[5];
// 对变量节点248传递过来的值进行组合
assign value_variable_to_check_124[35:30] = value_variable_248_to_check_124;
assign enable_variable_to_check_124[5] = enable_variable_248_to_check_124;


// 校验节点125的接口
wire [35:0] value_variable_to_check_125;
wire [35:0] value_check_125_to_variable;
wire [5:0] enable_variable_to_check_125;
wire [5:0] enable_check_125_to_variable;

// 拆分后校验节点125传递给变量节点6的值以及对变量节点6传递过来的值
wire [5:0] value_check_125_to_variable_6;
wire enable_check_125_to_variable_6;
wire [5:0] value_variable_6_to_check_125;
wire enable_variable_6_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_6 = value_check_125_to_variable[5:0];
assign enable_check_125_to_variable_6 = enable_check_125_to_variable[0];
// 对变量节点6传递过来的值进行组合
assign value_variable_to_check_125[5:0] = value_variable_6_to_check_125;
assign enable_variable_to_check_125[0] = enable_variable_6_to_check_125;

// 拆分后校验节点125传递给变量节点72的值以及对变量节点72传递过来的值
wire [5:0] value_check_125_to_variable_72;
wire enable_check_125_to_variable_72;
wire [5:0] value_variable_72_to_check_125;
wire enable_variable_72_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_72 = value_check_125_to_variable[11:6];
assign enable_check_125_to_variable_72 = enable_check_125_to_variable[1];
// 对变量节点72传递过来的值进行组合
assign value_variable_to_check_125[11:6] = value_variable_72_to_check_125;
assign enable_variable_to_check_125[1] = enable_variable_72_to_check_125;

// 拆分后校验节点125传递给变量节点126的值以及对变量节点126传递过来的值
wire [5:0] value_check_125_to_variable_126;
wire enable_check_125_to_variable_126;
wire [5:0] value_variable_126_to_check_125;
wire enable_variable_126_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_126 = value_check_125_to_variable[17:12];
assign enable_check_125_to_variable_126 = enable_check_125_to_variable[2];
// 对变量节点126传递过来的值进行组合
assign value_variable_to_check_125[17:12] = value_variable_126_to_check_125;
assign enable_variable_to_check_125[2] = enable_variable_126_to_check_125;

// 拆分后校验节点125传递给变量节点171的值以及对变量节点171传递过来的值
wire [5:0] value_check_125_to_variable_171;
wire enable_check_125_to_variable_171;
wire [5:0] value_variable_171_to_check_125;
wire enable_variable_171_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_171 = value_check_125_to_variable[23:18];
assign enable_check_125_to_variable_171 = enable_check_125_to_variable[3];
// 对变量节点171传递过来的值进行组合
assign value_variable_to_check_125[23:18] = value_variable_171_to_check_125;
assign enable_variable_to_check_125[3] = enable_variable_171_to_check_125;

// 拆分后校验节点125传递给变量节点212的值以及对变量节点212传递过来的值
wire [5:0] value_check_125_to_variable_212;
wire enable_check_125_to_variable_212;
wire [5:0] value_variable_212_to_check_125;
wire enable_variable_212_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_212 = value_check_125_to_variable[29:24];
assign enable_check_125_to_variable_212 = enable_check_125_to_variable[4];
// 对变量节点212传递过来的值进行组合
assign value_variable_to_check_125[29:24] = value_variable_212_to_check_125;
assign enable_variable_to_check_125[4] = enable_variable_212_to_check_125;

// 拆分后校验节点125传递给变量节点235的值以及对变量节点235传递过来的值
wire [5:0] value_check_125_to_variable_235;
wire enable_check_125_to_variable_235;
wire [5:0] value_variable_235_to_check_125;
wire enable_variable_235_to_check_125;
// 对校验节点125的输出值进行拆分
assign value_check_125_to_variable_235 = value_check_125_to_variable[35:30];
assign enable_check_125_to_variable_235 = enable_check_125_to_variable[5];
// 对变量节点235传递过来的值进行组合
assign value_variable_to_check_125[35:30] = value_variable_235_to_check_125;
assign enable_variable_to_check_125[5] = enable_variable_235_to_check_125;


// 校验节点126的接口
wire [35:0] value_variable_to_check_126;
wire [35:0] value_check_126_to_variable;
wire [5:0] enable_variable_to_check_126;
wire [5:0] enable_check_126_to_variable;

// 拆分后校验节点126传递给变量节点36的值以及对变量节点36传递过来的值
wire [5:0] value_check_126_to_variable_36;
wire enable_check_126_to_variable_36;
wire [5:0] value_variable_36_to_check_126;
wire enable_variable_36_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_36 = value_check_126_to_variable[5:0];
assign enable_check_126_to_variable_36 = enable_check_126_to_variable[0];
// 对变量节点36传递过来的值进行组合
assign value_variable_to_check_126[5:0] = value_variable_36_to_check_126;
assign enable_variable_to_check_126[0] = enable_variable_36_to_check_126;

// 拆分后校验节点126传递给变量节点76的值以及对变量节点76传递过来的值
wire [5:0] value_check_126_to_variable_76;
wire enable_check_126_to_variable_76;
wire [5:0] value_variable_76_to_check_126;
wire enable_variable_76_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_76 = value_check_126_to_variable[11:6];
assign enable_check_126_to_variable_76 = enable_check_126_to_variable[1];
// 对变量节点76传递过来的值进行组合
assign value_variable_to_check_126[11:6] = value_variable_76_to_check_126;
assign enable_variable_to_check_126[1] = enable_variable_76_to_check_126;

// 拆分后校验节点126传递给变量节点97的值以及对变量节点97传递过来的值
wire [5:0] value_check_126_to_variable_97;
wire enable_check_126_to_variable_97;
wire [5:0] value_variable_97_to_check_126;
wire enable_variable_97_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_97 = value_check_126_to_variable[17:12];
assign enable_check_126_to_variable_97 = enable_check_126_to_variable[2];
// 对变量节点97传递过来的值进行组合
assign value_variable_to_check_126[17:12] = value_variable_97_to_check_126;
assign enable_variable_to_check_126[2] = enable_variable_97_to_check_126;

// 拆分后校验节点126传递给变量节点154的值以及对变量节点154传递过来的值
wire [5:0] value_check_126_to_variable_154;
wire enable_check_126_to_variable_154;
wire [5:0] value_variable_154_to_check_126;
wire enable_variable_154_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_154 = value_check_126_to_variable[23:18];
assign enable_check_126_to_variable_154 = enable_check_126_to_variable[3];
// 对变量节点154传递过来的值进行组合
assign value_variable_to_check_126[23:18] = value_variable_154_to_check_126;
assign enable_variable_to_check_126[3] = enable_variable_154_to_check_126;

// 拆分后校验节点126传递给变量节点175的值以及对变量节点175传递过来的值
wire [5:0] value_check_126_to_variable_175;
wire enable_check_126_to_variable_175;
wire [5:0] value_variable_175_to_check_126;
wire enable_variable_175_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_175 = value_check_126_to_variable[29:24];
assign enable_check_126_to_variable_175 = enable_check_126_to_variable[4];
// 对变量节点175传递过来的值进行组合
assign value_variable_to_check_126[29:24] = value_variable_175_to_check_126;
assign enable_variable_to_check_126[4] = enable_variable_175_to_check_126;

// 拆分后校验节点126传递给变量节点244的值以及对变量节点244传递过来的值
wire [5:0] value_check_126_to_variable_244;
wire enable_check_126_to_variable_244;
wire [5:0] value_variable_244_to_check_126;
wire enable_variable_244_to_check_126;
// 对校验节点126的输出值进行拆分
assign value_check_126_to_variable_244 = value_check_126_to_variable[35:30];
assign enable_check_126_to_variable_244 = enable_check_126_to_variable[5];
// 对变量节点244传递过来的值进行组合
assign value_variable_to_check_126[35:30] = value_variable_244_to_check_126;
assign enable_variable_to_check_126[5] = enable_variable_244_to_check_126;


// 校验节点127的接口
wire [35:0] value_variable_to_check_127;
wire [35:0] value_check_127_to_variable;
wire [5:0] enable_variable_to_check_127;
wire [5:0] enable_check_127_to_variable;

// 拆分后校验节点127传递给变量节点23的值以及对变量节点23传递过来的值
wire [5:0] value_check_127_to_variable_23;
wire enable_check_127_to_variable_23;
wire [5:0] value_variable_23_to_check_127;
wire enable_variable_23_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_23 = value_check_127_to_variable[5:0];
assign enable_check_127_to_variable_23 = enable_check_127_to_variable[0];
// 对变量节点23传递过来的值进行组合
assign value_variable_to_check_127[5:0] = value_variable_23_to_check_127;
assign enable_variable_to_check_127[0] = enable_variable_23_to_check_127;

// 拆分后校验节点127传递给变量节点85的值以及对变量节点85传递过来的值
wire [5:0] value_check_127_to_variable_85;
wire enable_check_127_to_variable_85;
wire [5:0] value_variable_85_to_check_127;
wire enable_variable_85_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_85 = value_check_127_to_variable[11:6];
assign enable_check_127_to_variable_85 = enable_check_127_to_variable[1];
// 对变量节点85传递过来的值进行组合
assign value_variable_to_check_127[11:6] = value_variable_85_to_check_127;
assign enable_variable_to_check_127[1] = enable_variable_85_to_check_127;

// 拆分后校验节点127传递给变量节点125的值以及对变量节点125传递过来的值
wire [5:0] value_check_127_to_variable_125;
wire enable_check_127_to_variable_125;
wire [5:0] value_variable_125_to_check_127;
wire enable_variable_125_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_125 = value_check_127_to_variable[17:12];
assign enable_check_127_to_variable_125 = enable_check_127_to_variable[2];
// 对变量节点125传递过来的值进行组合
assign value_variable_to_check_127[17:12] = value_variable_125_to_check_127;
assign enable_variable_to_check_127[2] = enable_variable_125_to_check_127;

// 拆分后校验节点127传递给变量节点171的值以及对变量节点171传递过来的值
wire [5:0] value_check_127_to_variable_171;
wire enable_check_127_to_variable_171;
wire [5:0] value_variable_171_to_check_127;
wire enable_variable_171_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_171 = value_check_127_to_variable[23:18];
assign enable_check_127_to_variable_171 = enable_check_127_to_variable[3];
// 对变量节点171传递过来的值进行组合
assign value_variable_to_check_127[23:18] = value_variable_171_to_check_127;
assign enable_variable_to_check_127[3] = enable_variable_171_to_check_127;

// 拆分后校验节点127传递给变量节点185的值以及对变量节点185传递过来的值
wire [5:0] value_check_127_to_variable_185;
wire enable_check_127_to_variable_185;
wire [5:0] value_variable_185_to_check_127;
wire enable_variable_185_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_185 = value_check_127_to_variable[29:24];
assign enable_check_127_to_variable_185 = enable_check_127_to_variable[4];
// 对变量节点185传递过来的值进行组合
assign value_variable_to_check_127[29:24] = value_variable_185_to_check_127;
assign enable_variable_to_check_127[4] = enable_variable_185_to_check_127;

// 拆分后校验节点127传递给变量节点254的值以及对变量节点254传递过来的值
wire [5:0] value_check_127_to_variable_254;
wire enable_check_127_to_variable_254;
wire [5:0] value_variable_254_to_check_127;
wire enable_variable_254_to_check_127;
// 对校验节点127的输出值进行拆分
assign value_check_127_to_variable_254 = value_check_127_to_variable[35:30];
assign enable_check_127_to_variable_254 = enable_check_127_to_variable[5];
// 对变量节点254传递过来的值进行组合
assign value_variable_to_check_127[35:30] = value_variable_254_to_check_127;
assign enable_variable_to_check_127[5] = enable_variable_254_to_check_127;


// 变量节点0的接口
wire [17:0] value_check_to_variable_0;
wire [2:0] enable_check_to_variable_0;
wire [5:0] value_variable_0_to_decision;
wire [17:0] value_variable_0_to_check;

wire enable_variable_0_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_0[5:0] = value_check_0_to_variable_0;
assign enable_check_to_variable_0[0] = enable_check_0_to_variable_0;
// 将变量节点0的输出与校验节点0的输入相连
assign value_variable_0_to_check_0 = value_variable_0_to_check[5:0];
assign enable_variable_0_to_check_0 = enable_variable_0_to_check;

// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_0[11:6] = value_check_35_to_variable_0;
assign enable_check_to_variable_0[1] = enable_check_35_to_variable_0;
// 将变量节点0的输出与校验节点35的输入相连
assign value_variable_0_to_check_35 = value_variable_0_to_check[11:6];
assign enable_variable_0_to_check_35 = enable_variable_0_to_check;

// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_0[17:12] = value_check_100_to_variable_0;
assign enable_check_to_variable_0[2] = enable_check_100_to_variable_0;
// 将变量节点0的输出与校验节点100的输入相连
assign value_variable_0_to_check_100 = value_variable_0_to_check[17:12];
assign enable_variable_0_to_check_100 = enable_variable_0_to_check;


// 变量节点1的接口
wire [17:0] value_check_to_variable_1;
wire [2:0] enable_check_to_variable_1;
wire [5:0] value_variable_1_to_decision;
wire [17:0] value_variable_1_to_check;

wire enable_variable_1_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_1[5:0] = value_check_1_to_variable_1;
assign enable_check_to_variable_1[0] = enable_check_1_to_variable_1;
// 将变量节点1的输出与校验节点1的输入相连
assign value_variable_1_to_check_1 = value_variable_1_to_check[5:0];
assign enable_variable_1_to_check_1 = enable_variable_1_to_check;

// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_1[11:6] = value_check_6_to_variable_1;
assign enable_check_to_variable_1[1] = enable_check_6_to_variable_1;
// 将变量节点1的输出与校验节点6的输入相连
assign value_variable_1_to_check_6 = value_variable_1_to_check[11:6];
assign enable_variable_1_to_check_6 = enable_variable_1_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_1[17:12] = value_check_106_to_variable_1;
assign enable_check_to_variable_1[2] = enable_check_106_to_variable_1;
// 将变量节点1的输出与校验节点106的输入相连
assign value_variable_1_to_check_106 = value_variable_1_to_check[17:12];
assign enable_variable_1_to_check_106 = enable_variable_1_to_check;


// 变量节点2的接口
wire [17:0] value_check_to_variable_2;
wire [2:0] enable_check_to_variable_2;
wire [5:0] value_variable_2_to_decision;
wire [17:0] value_variable_2_to_check;

wire enable_variable_2_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_2[5:0] = value_check_2_to_variable_2;
assign enable_check_to_variable_2[0] = enable_check_2_to_variable_2;
// 将变量节点2的输出与校验节点2的输入相连
assign value_variable_2_to_check_2 = value_variable_2_to_check[5:0];
assign enable_variable_2_to_check_2 = enable_variable_2_to_check;

// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_2[11:6] = value_check_44_to_variable_2;
assign enable_check_to_variable_2[1] = enable_check_44_to_variable_2;
// 将变量节点2的输出与校验节点44的输入相连
assign value_variable_2_to_check_44 = value_variable_2_to_check[11:6];
assign enable_variable_2_to_check_44 = enable_variable_2_to_check;

// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_2[17:12] = value_check_99_to_variable_2;
assign enable_check_to_variable_2[2] = enable_check_99_to_variable_2;
// 将变量节点2的输出与校验节点99的输入相连
assign value_variable_2_to_check_99 = value_variable_2_to_check[17:12];
assign enable_variable_2_to_check_99 = enable_variable_2_to_check;


// 变量节点3的接口
wire [17:0] value_check_to_variable_3;
wire [2:0] enable_check_to_variable_3;
wire [5:0] value_variable_3_to_decision;
wire [17:0] value_variable_3_to_check;

wire enable_variable_3_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_3[5:0] = value_check_3_to_variable_3;
assign enable_check_to_variable_3[0] = enable_check_3_to_variable_3;
// 将变量节点3的输出与校验节点3的输入相连
assign value_variable_3_to_check_3 = value_variable_3_to_check[5:0];
assign enable_variable_3_to_check_3 = enable_variable_3_to_check;

// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_3[11:6] = value_check_74_to_variable_3;
assign enable_check_to_variable_3[1] = enable_check_74_to_variable_3;
// 将变量节点3的输出与校验节点74的输入相连
assign value_variable_3_to_check_74 = value_variable_3_to_check[11:6];
assign enable_variable_3_to_check_74 = enable_variable_3_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_3[17:12] = value_check_88_to_variable_3;
assign enable_check_to_variable_3[2] = enable_check_88_to_variable_3;
// 将变量节点3的输出与校验节点88的输入相连
assign value_variable_3_to_check_88 = value_variable_3_to_check[17:12];
assign enable_variable_3_to_check_88 = enable_variable_3_to_check;


// 变量节点4的接口
wire [17:0] value_check_to_variable_4;
wire [2:0] enable_check_to_variable_4;
wire [5:0] value_variable_4_to_decision;
wire [17:0] value_variable_4_to_check;

wire enable_variable_4_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_4[5:0] = value_check_4_to_variable_4;
assign enable_check_to_variable_4[0] = enable_check_4_to_variable_4;
// 将变量节点4的输出与校验节点4的输入相连
assign value_variable_4_to_check_4 = value_variable_4_to_check[5:0];
assign enable_variable_4_to_check_4 = enable_variable_4_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_4[11:6] = value_check_91_to_variable_4;
assign enable_check_to_variable_4[1] = enable_check_91_to_variable_4;
// 将变量节点4的输出与校验节点91的输入相连
assign value_variable_4_to_check_91 = value_variable_4_to_check[11:6];
assign enable_variable_4_to_check_91 = enable_variable_4_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_4[17:12] = value_check_101_to_variable_4;
assign enable_check_to_variable_4[2] = enable_check_101_to_variable_4;
// 将变量节点4的输出与校验节点101的输入相连
assign value_variable_4_to_check_101 = value_variable_4_to_check[17:12];
assign enable_variable_4_to_check_101 = enable_variable_4_to_check;


// 变量节点5的接口
wire [17:0] value_check_to_variable_5;
wire [2:0] enable_check_to_variable_5;
wire [5:0] value_variable_5_to_decision;
wire [17:0] value_variable_5_to_check;

wire enable_variable_5_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_5[5:0] = value_check_5_to_variable_5;
assign enable_check_to_variable_5[0] = enable_check_5_to_variable_5;
// 将变量节点5的输出与校验节点5的输入相连
assign value_variable_5_to_check_5 = value_variable_5_to_check[5:0];
assign enable_variable_5_to_check_5 = enable_variable_5_to_check;

// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_5[11:6] = value_check_46_to_variable_5;
assign enable_check_to_variable_5[1] = enable_check_46_to_variable_5;
// 将变量节点5的输出与校验节点46的输入相连
assign value_variable_5_to_check_46 = value_variable_5_to_check[11:6];
assign enable_variable_5_to_check_46 = enable_variable_5_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_5[17:12] = value_check_114_to_variable_5;
assign enable_check_to_variable_5[2] = enable_check_114_to_variable_5;
// 将变量节点5的输出与校验节点114的输入相连
assign value_variable_5_to_check_114 = value_variable_5_to_check[17:12];
assign enable_variable_5_to_check_114 = enable_variable_5_to_check;


// 变量节点6的接口
wire [17:0] value_check_to_variable_6;
wire [2:0] enable_check_to_variable_6;
wire [5:0] value_variable_6_to_decision;
wire [17:0] value_variable_6_to_check;

wire enable_variable_6_to_check;
// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_6[5:0] = value_check_7_to_variable_6;
assign enable_check_to_variable_6[0] = enable_check_7_to_variable_6;
// 将变量节点6的输出与校验节点7的输入相连
assign value_variable_6_to_check_7 = value_variable_6_to_check[5:0];
assign enable_variable_6_to_check_7 = enable_variable_6_to_check;

// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_6[11:6] = value_check_73_to_variable_6;
assign enable_check_to_variable_6[1] = enable_check_73_to_variable_6;
// 将变量节点6的输出与校验节点73的输入相连
assign value_variable_6_to_check_73 = value_variable_6_to_check[11:6];
assign enable_variable_6_to_check_73 = enable_variable_6_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_6[17:12] = value_check_125_to_variable_6;
assign enable_check_to_variable_6[2] = enable_check_125_to_variable_6;
// 将变量节点6的输出与校验节点125的输入相连
assign value_variable_6_to_check_125 = value_variable_6_to_check[17:12];
assign enable_variable_6_to_check_125 = enable_variable_6_to_check;


// 变量节点7的接口
wire [17:0] value_check_to_variable_7;
wire [2:0] enable_check_to_variable_7;
wire [5:0] value_variable_7_to_decision;
wire [17:0] value_variable_7_to_check;

wire enable_variable_7_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_7[5:0] = value_check_8_to_variable_7;
assign enable_check_to_variable_7[0] = enable_check_8_to_variable_7;
// 将变量节点7的输出与校验节点8的输入相连
assign value_variable_7_to_check_8 = value_variable_7_to_check[5:0];
assign enable_variable_7_to_check_8 = enable_variable_7_to_check;

// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_7[11:6] = value_check_51_to_variable_7;
assign enable_check_to_variable_7[1] = enable_check_51_to_variable_7;
// 将变量节点7的输出与校验节点51的输入相连
assign value_variable_7_to_check_51 = value_variable_7_to_check[11:6];
assign enable_variable_7_to_check_51 = enable_variable_7_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_7[17:12] = value_check_61_to_variable_7;
assign enable_check_to_variable_7[2] = enable_check_61_to_variable_7;
// 将变量节点7的输出与校验节点61的输入相连
assign value_variable_7_to_check_61 = value_variable_7_to_check[17:12];
assign enable_variable_7_to_check_61 = enable_variable_7_to_check;


// 变量节点8的接口
wire [17:0] value_check_to_variable_8;
wire [2:0] enable_check_to_variable_8;
wire [5:0] value_variable_8_to_decision;
wire [17:0] value_variable_8_to_check;

wire enable_variable_8_to_check;
// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_8[5:0] = value_check_9_to_variable_8;
assign enable_check_to_variable_8[0] = enable_check_9_to_variable_8;
// 将变量节点8的输出与校验节点9的输入相连
assign value_variable_8_to_check_9 = value_variable_8_to_check[5:0];
assign enable_variable_8_to_check_9 = enable_variable_8_to_check;

// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_8[11:6] = value_check_57_to_variable_8;
assign enable_check_to_variable_8[1] = enable_check_57_to_variable_8;
// 将变量节点8的输出与校验节点57的输入相连
assign value_variable_8_to_check_57 = value_variable_8_to_check[11:6];
assign enable_variable_8_to_check_57 = enable_variable_8_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_8[17:12] = value_check_93_to_variable_8;
assign enable_check_to_variable_8[2] = enable_check_93_to_variable_8;
// 将变量节点8的输出与校验节点93的输入相连
assign value_variable_8_to_check_93 = value_variable_8_to_check[17:12];
assign enable_variable_8_to_check_93 = enable_variable_8_to_check;


// 变量节点9的接口
wire [17:0] value_check_to_variable_9;
wire [2:0] enable_check_to_variable_9;
wire [5:0] value_variable_9_to_decision;
wire [17:0] value_variable_9_to_check;

wire enable_variable_9_to_check;
// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_9[5:0] = value_check_10_to_variable_9;
assign enable_check_to_variable_9[0] = enable_check_10_to_variable_9;
// 将变量节点9的输出与校验节点10的输入相连
assign value_variable_9_to_check_10 = value_variable_9_to_check[5:0];
assign enable_variable_9_to_check_10 = enable_variable_9_to_check;

// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_9[11:6] = value_check_14_to_variable_9;
assign enable_check_to_variable_9[1] = enable_check_14_to_variable_9;
// 将变量节点9的输出与校验节点14的输入相连
assign value_variable_9_to_check_14 = value_variable_9_to_check[11:6];
assign enable_variable_9_to_check_14 = enable_variable_9_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_9[17:12] = value_check_94_to_variable_9;
assign enable_check_to_variable_9[2] = enable_check_94_to_variable_9;
// 将变量节点9的输出与校验节点94的输入相连
assign value_variable_9_to_check_94 = value_variable_9_to_check[17:12];
assign enable_variable_9_to_check_94 = enable_variable_9_to_check;


// 变量节点10的接口
wire [17:0] value_check_to_variable_10;
wire [2:0] enable_check_to_variable_10;
wire [5:0] value_variable_10_to_decision;
wire [17:0] value_variable_10_to_check;

wire enable_variable_10_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_10[5:0] = value_check_11_to_variable_10;
assign enable_check_to_variable_10[0] = enable_check_11_to_variable_10;
// 将变量节点10的输出与校验节点11的输入相连
assign value_variable_10_to_check_11 = value_variable_10_to_check[5:0];
assign enable_variable_10_to_check_11 = enable_variable_10_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_10[11:6] = value_check_107_to_variable_10;
assign enable_check_to_variable_10[1] = enable_check_107_to_variable_10;
// 将变量节点10的输出与校验节点107的输入相连
assign value_variable_10_to_check_107 = value_variable_10_to_check[11:6];
assign enable_variable_10_to_check_107 = enable_variable_10_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_10[17:12] = value_check_111_to_variable_10;
assign enable_check_to_variable_10[2] = enable_check_111_to_variable_10;
// 将变量节点10的输出与校验节点111的输入相连
assign value_variable_10_to_check_111 = value_variable_10_to_check[17:12];
assign enable_variable_10_to_check_111 = enable_variable_10_to_check;


// 变量节点11的接口
wire [17:0] value_check_to_variable_11;
wire [2:0] enable_check_to_variable_11;
wire [5:0] value_variable_11_to_decision;
wire [17:0] value_variable_11_to_check;

wire enable_variable_11_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_11[5:0] = value_check_12_to_variable_11;
assign enable_check_to_variable_11[0] = enable_check_12_to_variable_11;
// 将变量节点11的输出与校验节点12的输入相连
assign value_variable_11_to_check_12 = value_variable_11_to_check[5:0];
assign enable_variable_11_to_check_12 = enable_variable_11_to_check;

// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_11[11:6] = value_check_29_to_variable_11;
assign enable_check_to_variable_11[1] = enable_check_29_to_variable_11;
// 将变量节点11的输出与校验节点29的输入相连
assign value_variable_11_to_check_29 = value_variable_11_to_check[11:6];
assign enable_variable_11_to_check_29 = enable_variable_11_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_11[17:12] = value_check_117_to_variable_11;
assign enable_check_to_variable_11[2] = enable_check_117_to_variable_11;
// 将变量节点11的输出与校验节点117的输入相连
assign value_variable_11_to_check_117 = value_variable_11_to_check[17:12];
assign enable_variable_11_to_check_117 = enable_variable_11_to_check;


// 变量节点12的接口
wire [17:0] value_check_to_variable_12;
wire [2:0] enable_check_to_variable_12;
wire [5:0] value_variable_12_to_decision;
wire [17:0] value_variable_12_to_check;

wire enable_variable_12_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_12[5:0] = value_check_13_to_variable_12;
assign enable_check_to_variable_12[0] = enable_check_13_to_variable_12;
// 将变量节点12的输出与校验节点13的输入相连
assign value_variable_12_to_check_13 = value_variable_12_to_check[5:0];
assign enable_variable_12_to_check_13 = enable_variable_12_to_check;

// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_12[11:6] = value_check_15_to_variable_12;
assign enable_check_to_variable_12[1] = enable_check_15_to_variable_12;
// 将变量节点12的输出与校验节点15的输入相连
assign value_variable_12_to_check_15 = value_variable_12_to_check[11:6];
assign enable_variable_12_to_check_15 = enable_variable_12_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_12[17:12] = value_check_119_to_variable_12;
assign enable_check_to_variable_12[2] = enable_check_119_to_variable_12;
// 将变量节点12的输出与校验节点119的输入相连
assign value_variable_12_to_check_119 = value_variable_12_to_check[17:12];
assign enable_variable_12_to_check_119 = enable_variable_12_to_check;


// 变量节点13的接口
wire [17:0] value_check_to_variable_13;
wire [2:0] enable_check_to_variable_13;
wire [5:0] value_variable_13_to_decision;
wire [17:0] value_variable_13_to_check;

wire enable_variable_13_to_check;
// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_13[5:0] = value_check_16_to_variable_13;
assign enable_check_to_variable_13[0] = enable_check_16_to_variable_13;
// 将变量节点13的输出与校验节点16的输入相连
assign value_variable_13_to_check_16 = value_variable_13_to_check[5:0];
assign enable_variable_13_to_check_16 = enable_variable_13_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_13[11:6] = value_check_81_to_variable_13;
assign enable_check_to_variable_13[1] = enable_check_81_to_variable_13;
// 将变量节点13的输出与校验节点81的输入相连
assign value_variable_13_to_check_81 = value_variable_13_to_check[11:6];
assign enable_variable_13_to_check_81 = enable_variable_13_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_13[17:12] = value_check_96_to_variable_13;
assign enable_check_to_variable_13[2] = enable_check_96_to_variable_13;
// 将变量节点13的输出与校验节点96的输入相连
assign value_variable_13_to_check_96 = value_variable_13_to_check[17:12];
assign enable_variable_13_to_check_96 = enable_variable_13_to_check;


// 变量节点14的接口
wire [17:0] value_check_to_variable_14;
wire [2:0] enable_check_to_variable_14;
wire [5:0] value_variable_14_to_decision;
wire [17:0] value_variable_14_to_check;

wire enable_variable_14_to_check;
// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_14[5:0] = value_check_17_to_variable_14;
assign enable_check_to_variable_14[0] = enable_check_17_to_variable_14;
// 将变量节点14的输出与校验节点17的输入相连
assign value_variable_14_to_check_17 = value_variable_14_to_check[5:0];
assign enable_variable_14_to_check_17 = enable_variable_14_to_check;

// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_14[11:6] = value_check_76_to_variable_14;
assign enable_check_to_variable_14[1] = enable_check_76_to_variable_14;
// 将变量节点14的输出与校验节点76的输入相连
assign value_variable_14_to_check_76 = value_variable_14_to_check[11:6];
assign enable_variable_14_to_check_76 = enable_variable_14_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_14[17:12] = value_check_90_to_variable_14;
assign enable_check_to_variable_14[2] = enable_check_90_to_variable_14;
// 将变量节点14的输出与校验节点90的输入相连
assign value_variable_14_to_check_90 = value_variable_14_to_check[17:12];
assign enable_variable_14_to_check_90 = enable_variable_14_to_check;


// 变量节点15的接口
wire [17:0] value_check_to_variable_15;
wire [2:0] enable_check_to_variable_15;
wire [5:0] value_variable_15_to_decision;
wire [17:0] value_variable_15_to_check;

wire enable_variable_15_to_check;
// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_15[5:0] = value_check_18_to_variable_15;
assign enable_check_to_variable_15[0] = enable_check_18_to_variable_15;
// 将变量节点15的输出与校验节点18的输入相连
assign value_variable_15_to_check_18 = value_variable_15_to_check[5:0];
assign enable_variable_15_to_check_18 = enable_variable_15_to_check;

// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_15[11:6] = value_check_40_to_variable_15;
assign enable_check_to_variable_15[1] = enable_check_40_to_variable_15;
// 将变量节点15的输出与校验节点40的输入相连
assign value_variable_15_to_check_40 = value_variable_15_to_check[11:6];
assign enable_variable_15_to_check_40 = enable_variable_15_to_check;

// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_15[17:12] = value_check_72_to_variable_15;
assign enable_check_to_variable_15[2] = enable_check_72_to_variable_15;
// 将变量节点15的输出与校验节点72的输入相连
assign value_variable_15_to_check_72 = value_variable_15_to_check[17:12];
assign enable_variable_15_to_check_72 = enable_variable_15_to_check;


// 变量节点16的接口
wire [17:0] value_check_to_variable_16;
wire [2:0] enable_check_to_variable_16;
wire [5:0] value_variable_16_to_decision;
wire [17:0] value_variable_16_to_check;

wire enable_variable_16_to_check;
// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_16[5:0] = value_check_19_to_variable_16;
assign enable_check_to_variable_16[0] = enable_check_19_to_variable_16;
// 将变量节点16的输出与校验节点19的输入相连
assign value_variable_16_to_check_19 = value_variable_16_to_check[5:0];
assign enable_variable_16_to_check_19 = enable_variable_16_to_check;

// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_16[11:6] = value_check_95_to_variable_16;
assign enable_check_to_variable_16[1] = enable_check_95_to_variable_16;
// 将变量节点16的输出与校验节点95的输入相连
assign value_variable_16_to_check_95 = value_variable_16_to_check[11:6];
assign enable_variable_16_to_check_95 = enable_variable_16_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_16[17:12] = value_check_121_to_variable_16;
assign enable_check_to_variable_16[2] = enable_check_121_to_variable_16;
// 将变量节点16的输出与校验节点121的输入相连
assign value_variable_16_to_check_121 = value_variable_16_to_check[17:12];
assign enable_variable_16_to_check_121 = enable_variable_16_to_check;


// 变量节点17的接口
wire [17:0] value_check_to_variable_17;
wire [2:0] enable_check_to_variable_17;
wire [5:0] value_variable_17_to_decision;
wire [17:0] value_variable_17_to_check;

wire enable_variable_17_to_check;
// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_17[5:0] = value_check_20_to_variable_17;
assign enable_check_to_variable_17[0] = enable_check_20_to_variable_17;
// 将变量节点17的输出与校验节点20的输入相连
assign value_variable_17_to_check_20 = value_variable_17_to_check[5:0];
assign enable_variable_17_to_check_20 = enable_variable_17_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_17[11:6] = value_check_34_to_variable_17;
assign enable_check_to_variable_17[1] = enable_check_34_to_variable_17;
// 将变量节点17的输出与校验节点34的输入相连
assign value_variable_17_to_check_34 = value_variable_17_to_check[11:6];
assign enable_variable_17_to_check_34 = enable_variable_17_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_17[17:12] = value_check_104_to_variable_17;
assign enable_check_to_variable_17[2] = enable_check_104_to_variable_17;
// 将变量节点17的输出与校验节点104的输入相连
assign value_variable_17_to_check_104 = value_variable_17_to_check[17:12];
assign enable_variable_17_to_check_104 = enable_variable_17_to_check;


// 变量节点18的接口
wire [17:0] value_check_to_variable_18;
wire [2:0] enable_check_to_variable_18;
wire [5:0] value_variable_18_to_decision;
wire [17:0] value_variable_18_to_check;

wire enable_variable_18_to_check;
// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_18[5:0] = value_check_21_to_variable_18;
assign enable_check_to_variable_18[0] = enable_check_21_to_variable_18;
// 将变量节点18的输出与校验节点21的输入相连
assign value_variable_18_to_check_21 = value_variable_18_to_check[5:0];
assign enable_variable_18_to_check_21 = enable_variable_18_to_check;

// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_18[11:6] = value_check_22_to_variable_18;
assign enable_check_to_variable_18[1] = enable_check_22_to_variable_18;
// 将变量节点18的输出与校验节点22的输入相连
assign value_variable_18_to_check_22 = value_variable_18_to_check[11:6];
assign enable_variable_18_to_check_22 = enable_variable_18_to_check;

// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_18[17:12] = value_check_56_to_variable_18;
assign enable_check_to_variable_18[2] = enable_check_56_to_variable_18;
// 将变量节点18的输出与校验节点56的输入相连
assign value_variable_18_to_check_56 = value_variable_18_to_check[17:12];
assign enable_variable_18_to_check_56 = enable_variable_18_to_check;


// 变量节点19的接口
wire [17:0] value_check_to_variable_19;
wire [2:0] enable_check_to_variable_19;
wire [5:0] value_variable_19_to_decision;
wire [17:0] value_variable_19_to_check;

wire enable_variable_19_to_check;
// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_19[5:0] = value_check_23_to_variable_19;
assign enable_check_to_variable_19[0] = enable_check_23_to_variable_19;
// 将变量节点19的输出与校验节点23的输入相连
assign value_variable_19_to_check_23 = value_variable_19_to_check[5:0];
assign enable_variable_19_to_check_23 = enable_variable_19_to_check;

// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_19[11:6] = value_check_37_to_variable_19;
assign enable_check_to_variable_19[1] = enable_check_37_to_variable_19;
// 将变量节点19的输出与校验节点37的输入相连
assign value_variable_19_to_check_37 = value_variable_19_to_check[11:6];
assign enable_variable_19_to_check_37 = enable_variable_19_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_19[17:12] = value_check_105_to_variable_19;
assign enable_check_to_variable_19[2] = enable_check_105_to_variable_19;
// 将变量节点19的输出与校验节点105的输入相连
assign value_variable_19_to_check_105 = value_variable_19_to_check[17:12];
assign enable_variable_19_to_check_105 = enable_variable_19_to_check;


// 变量节点20的接口
wire [17:0] value_check_to_variable_20;
wire [2:0] enable_check_to_variable_20;
wire [5:0] value_variable_20_to_decision;
wire [17:0] value_variable_20_to_check;

wire enable_variable_20_to_check;
// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_20[5:0] = value_check_24_to_variable_20;
assign enable_check_to_variable_20[0] = enable_check_24_to_variable_20;
// 将变量节点20的输出与校验节点24的输入相连
assign value_variable_20_to_check_24 = value_variable_20_to_check[5:0];
assign enable_variable_20_to_check_24 = enable_variable_20_to_check;

// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_20[11:6] = value_check_36_to_variable_20;
assign enable_check_to_variable_20[1] = enable_check_36_to_variable_20;
// 将变量节点20的输出与校验节点36的输入相连
assign value_variable_20_to_check_36 = value_variable_20_to_check[11:6];
assign enable_variable_20_to_check_36 = enable_variable_20_to_check;

// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_20[17:12] = value_check_41_to_variable_20;
assign enable_check_to_variable_20[2] = enable_check_41_to_variable_20;
// 将变量节点20的输出与校验节点41的输入相连
assign value_variable_20_to_check_41 = value_variable_20_to_check[17:12];
assign enable_variable_20_to_check_41 = enable_variable_20_to_check;


// 变量节点21的接口
wire [17:0] value_check_to_variable_21;
wire [2:0] enable_check_to_variable_21;
wire [5:0] value_variable_21_to_decision;
wire [17:0] value_variable_21_to_check;

wire enable_variable_21_to_check;
// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_21[5:0] = value_check_25_to_variable_21;
assign enable_check_to_variable_21[0] = enable_check_25_to_variable_21;
// 将变量节点21的输出与校验节点25的输入相连
assign value_variable_21_to_check_25 = value_variable_21_to_check[5:0];
assign enable_variable_21_to_check_25 = enable_variable_21_to_check;

// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_21[11:6] = value_check_39_to_variable_21;
assign enable_check_to_variable_21[1] = enable_check_39_to_variable_21;
// 将变量节点21的输出与校验节点39的输入相连
assign value_variable_21_to_check_39 = value_variable_21_to_check[11:6];
assign enable_variable_21_to_check_39 = enable_variable_21_to_check;

// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_21[17:12] = value_check_48_to_variable_21;
assign enable_check_to_variable_21[2] = enable_check_48_to_variable_21;
// 将变量节点21的输出与校验节点48的输入相连
assign value_variable_21_to_check_48 = value_variable_21_to_check[17:12];
assign enable_variable_21_to_check_48 = enable_variable_21_to_check;


// 变量节点22的接口
wire [17:0] value_check_to_variable_22;
wire [2:0] enable_check_to_variable_22;
wire [5:0] value_variable_22_to_decision;
wire [17:0] value_variable_22_to_check;

wire enable_variable_22_to_check;
// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_22[5:0] = value_check_26_to_variable_22;
assign enable_check_to_variable_22[0] = enable_check_26_to_variable_22;
// 将变量节点22的输出与校验节点26的输入相连
assign value_variable_22_to_check_26 = value_variable_22_to_check[5:0];
assign enable_variable_22_to_check_26 = enable_variable_22_to_check;

// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_22[11:6] = value_check_63_to_variable_22;
assign enable_check_to_variable_22[1] = enable_check_63_to_variable_22;
// 将变量节点22的输出与校验节点63的输入相连
assign value_variable_22_to_check_63 = value_variable_22_to_check[11:6];
assign enable_variable_22_to_check_63 = enable_variable_22_to_check;

// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_22[17:12] = value_check_66_to_variable_22;
assign enable_check_to_variable_22[2] = enable_check_66_to_variable_22;
// 将变量节点22的输出与校验节点66的输入相连
assign value_variable_22_to_check_66 = value_variable_22_to_check[17:12];
assign enable_variable_22_to_check_66 = enable_variable_22_to_check;


// 变量节点23的接口
wire [17:0] value_check_to_variable_23;
wire [2:0] enable_check_to_variable_23;
wire [5:0] value_variable_23_to_decision;
wire [17:0] value_variable_23_to_check;

wire enable_variable_23_to_check;
// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_23[5:0] = value_check_27_to_variable_23;
assign enable_check_to_variable_23[0] = enable_check_27_to_variable_23;
// 将变量节点23的输出与校验节点27的输入相连
assign value_variable_23_to_check_27 = value_variable_23_to_check[5:0];
assign enable_variable_23_to_check_27 = enable_variable_23_to_check;

// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_23[11:6] = value_check_62_to_variable_23;
assign enable_check_to_variable_23[1] = enable_check_62_to_variable_23;
// 将变量节点23的输出与校验节点62的输入相连
assign value_variable_23_to_check_62 = value_variable_23_to_check[11:6];
assign enable_variable_23_to_check_62 = enable_variable_23_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_23[17:12] = value_check_127_to_variable_23;
assign enable_check_to_variable_23[2] = enable_check_127_to_variable_23;
// 将变量节点23的输出与校验节点127的输入相连
assign value_variable_23_to_check_127 = value_variable_23_to_check[17:12];
assign enable_variable_23_to_check_127 = enable_variable_23_to_check;


// 变量节点24的接口
wire [17:0] value_check_to_variable_24;
wire [2:0] enable_check_to_variable_24;
wire [5:0] value_variable_24_to_decision;
wire [17:0] value_variable_24_to_check;

wire enable_variable_24_to_check;
// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_24[5:0] = value_check_28_to_variable_24;
assign enable_check_to_variable_24[0] = enable_check_28_to_variable_24;
// 将变量节点24的输出与校验节点28的输入相连
assign value_variable_24_to_check_28 = value_variable_24_to_check[5:0];
assign enable_variable_24_to_check_28 = enable_variable_24_to_check;

// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_24[11:6] = value_check_59_to_variable_24;
assign enable_check_to_variable_24[1] = enable_check_59_to_variable_24;
// 将变量节点24的输出与校验节点59的输入相连
assign value_variable_24_to_check_59 = value_variable_24_to_check[11:6];
assign enable_variable_24_to_check_59 = enable_variable_24_to_check;

// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_24[17:12] = value_check_65_to_variable_24;
assign enable_check_to_variable_24[2] = enable_check_65_to_variable_24;
// 将变量节点24的输出与校验节点65的输入相连
assign value_variable_24_to_check_65 = value_variable_24_to_check[17:12];
assign enable_variable_24_to_check_65 = enable_variable_24_to_check;


// 变量节点25的接口
wire [17:0] value_check_to_variable_25;
wire [2:0] enable_check_to_variable_25;
wire [5:0] value_variable_25_to_decision;
wire [17:0] value_variable_25_to_check;

wire enable_variable_25_to_check;
// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_25[5:0] = value_check_30_to_variable_25;
assign enable_check_to_variable_25[0] = enable_check_30_to_variable_25;
// 将变量节点25的输出与校验节点30的输入相连
assign value_variable_25_to_check_30 = value_variable_25_to_check[5:0];
assign enable_variable_25_to_check_30 = enable_variable_25_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_25[11:6] = value_check_85_to_variable_25;
assign enable_check_to_variable_25[1] = enable_check_85_to_variable_25;
// 将变量节点25的输出与校验节点85的输入相连
assign value_variable_25_to_check_85 = value_variable_25_to_check[11:6];
assign enable_variable_25_to_check_85 = enable_variable_25_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_25[17:12] = value_check_116_to_variable_25;
assign enable_check_to_variable_25[2] = enable_check_116_to_variable_25;
// 将变量节点25的输出与校验节点116的输入相连
assign value_variable_25_to_check_116 = value_variable_25_to_check[17:12];
assign enable_variable_25_to_check_116 = enable_variable_25_to_check;


// 变量节点26的接口
wire [17:0] value_check_to_variable_26;
wire [2:0] enable_check_to_variable_26;
wire [5:0] value_variable_26_to_decision;
wire [17:0] value_variable_26_to_check;

wire enable_variable_26_to_check;
// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_26[5:0] = value_check_31_to_variable_26;
assign enable_check_to_variable_26[0] = enable_check_31_to_variable_26;
// 将变量节点26的输出与校验节点31的输入相连
assign value_variable_26_to_check_31 = value_variable_26_to_check[5:0];
assign enable_variable_26_to_check_31 = enable_variable_26_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_26[11:6] = value_check_75_to_variable_26;
assign enable_check_to_variable_26[1] = enable_check_75_to_variable_26;
// 将变量节点26的输出与校验节点75的输入相连
assign value_variable_26_to_check_75 = value_variable_26_to_check[11:6];
assign enable_variable_26_to_check_75 = enable_variable_26_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_26[17:12] = value_check_113_to_variable_26;
assign enable_check_to_variable_26[2] = enable_check_113_to_variable_26;
// 将变量节点26的输出与校验节点113的输入相连
assign value_variable_26_to_check_113 = value_variable_26_to_check[17:12];
assign enable_variable_26_to_check_113 = enable_variable_26_to_check;


// 变量节点27的接口
wire [17:0] value_check_to_variable_27;
wire [2:0] enable_check_to_variable_27;
wire [5:0] value_variable_27_to_decision;
wire [17:0] value_variable_27_to_check;

wire enable_variable_27_to_check;
// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_27[5:0] = value_check_32_to_variable_27;
assign enable_check_to_variable_27[0] = enable_check_32_to_variable_27;
// 将变量节点27的输出与校验节点32的输入相连
assign value_variable_27_to_check_32 = value_variable_27_to_check[5:0];
assign enable_variable_27_to_check_32 = enable_variable_27_to_check;

// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_27[11:6] = value_check_38_to_variable_27;
assign enable_check_to_variable_27[1] = enable_check_38_to_variable_27;
// 将变量节点27的输出与校验节点38的输入相连
assign value_variable_27_to_check_38 = value_variable_27_to_check[11:6];
assign enable_variable_27_to_check_38 = enable_variable_27_to_check;

// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_27[17:12] = value_check_110_to_variable_27;
assign enable_check_to_variable_27[2] = enable_check_110_to_variable_27;
// 将变量节点27的输出与校验节点110的输入相连
assign value_variable_27_to_check_110 = value_variable_27_to_check[17:12];
assign enable_variable_27_to_check_110 = enable_variable_27_to_check;


// 变量节点28的接口
wire [17:0] value_check_to_variable_28;
wire [2:0] enable_check_to_variable_28;
wire [5:0] value_variable_28_to_decision;
wire [17:0] value_variable_28_to_check;

wire enable_variable_28_to_check;
// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_28[5:0] = value_check_33_to_variable_28;
assign enable_check_to_variable_28[0] = enable_check_33_to_variable_28;
// 将变量节点28的输出与校验节点33的输入相连
assign value_variable_28_to_check_33 = value_variable_28_to_check[5:0];
assign enable_variable_28_to_check_33 = enable_variable_28_to_check;

// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_28[11:6] = value_check_42_to_variable_28;
assign enable_check_to_variable_28[1] = enable_check_42_to_variable_28;
// 将变量节点28的输出与校验节点42的输入相连
assign value_variable_28_to_check_42 = value_variable_28_to_check[11:6];
assign enable_variable_28_to_check_42 = enable_variable_28_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_28[17:12] = value_check_84_to_variable_28;
assign enable_check_to_variable_28[2] = enable_check_84_to_variable_28;
// 将变量节点28的输出与校验节点84的输入相连
assign value_variable_28_to_check_84 = value_variable_28_to_check[17:12];
assign enable_variable_28_to_check_84 = enable_variable_28_to_check;


// 变量节点29的接口
wire [17:0] value_check_to_variable_29;
wire [2:0] enable_check_to_variable_29;
wire [5:0] value_variable_29_to_decision;
wire [17:0] value_variable_29_to_check;

wire enable_variable_29_to_check;
// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_29[5:0] = value_check_43_to_variable_29;
assign enable_check_to_variable_29[0] = enable_check_43_to_variable_29;
// 将变量节点29的输出与校验节点43的输入相连
assign value_variable_29_to_check_43 = value_variable_29_to_check[5:0];
assign enable_variable_29_to_check_43 = enable_variable_29_to_check;

// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_29[11:6] = value_check_83_to_variable_29;
assign enable_check_to_variable_29[1] = enable_check_83_to_variable_29;
// 将变量节点29的输出与校验节点83的输入相连
assign value_variable_29_to_check_83 = value_variable_29_to_check[11:6];
assign enable_variable_29_to_check_83 = enable_variable_29_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_29[17:12] = value_check_87_to_variable_29;
assign enable_check_to_variable_29[2] = enable_check_87_to_variable_29;
// 将变量节点29的输出与校验节点87的输入相连
assign value_variable_29_to_check_87 = value_variable_29_to_check[17:12];
assign enable_variable_29_to_check_87 = enable_variable_29_to_check;


// 变量节点30的接口
wire [17:0] value_check_to_variable_30;
wire [2:0] enable_check_to_variable_30;
wire [5:0] value_variable_30_to_decision;
wire [17:0] value_variable_30_to_check;

wire enable_variable_30_to_check;
// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_30[5:0] = value_check_45_to_variable_30;
assign enable_check_to_variable_30[0] = enable_check_45_to_variable_30;
// 将变量节点30的输出与校验节点45的输入相连
assign value_variable_30_to_check_45 = value_variable_30_to_check[5:0];
assign enable_variable_30_to_check_45 = enable_variable_30_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_30[11:6] = value_check_120_to_variable_30;
assign enable_check_to_variable_30[1] = enable_check_120_to_variable_30;
// 将变量节点30的输出与校验节点120的输入相连
assign value_variable_30_to_check_120 = value_variable_30_to_check[11:6];
assign enable_variable_30_to_check_120 = enable_variable_30_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_30[17:12] = value_check_124_to_variable_30;
assign enable_check_to_variable_30[2] = enable_check_124_to_variable_30;
// 将变量节点30的输出与校验节点124的输入相连
assign value_variable_30_to_check_124 = value_variable_30_to_check[17:12];
assign enable_variable_30_to_check_124 = enable_variable_30_to_check;


// 变量节点31的接口
wire [17:0] value_check_to_variable_31;
wire [2:0] enable_check_to_variable_31;
wire [5:0] value_variable_31_to_decision;
wire [17:0] value_variable_31_to_check;

wire enable_variable_31_to_check;
// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_31[5:0] = value_check_47_to_variable_31;
assign enable_check_to_variable_31[0] = enable_check_47_to_variable_31;
// 将变量节点31的输出与校验节点47的输入相连
assign value_variable_31_to_check_47 = value_variable_31_to_check[5:0];
assign enable_variable_31_to_check_47 = enable_variable_31_to_check;

// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_31[11:6] = value_check_54_to_variable_31;
assign enable_check_to_variable_31[1] = enable_check_54_to_variable_31;
// 将变量节点31的输出与校验节点54的输入相连
assign value_variable_31_to_check_54 = value_variable_31_to_check[11:6];
assign enable_variable_31_to_check_54 = enable_variable_31_to_check;

// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_31[17:12] = value_check_67_to_variable_31;
assign enable_check_to_variable_31[2] = enable_check_67_to_variable_31;
// 将变量节点31的输出与校验节点67的输入相连
assign value_variable_31_to_check_67 = value_variable_31_to_check[17:12];
assign enable_variable_31_to_check_67 = enable_variable_31_to_check;


// 变量节点32的接口
wire [17:0] value_check_to_variable_32;
wire [2:0] enable_check_to_variable_32;
wire [5:0] value_variable_32_to_decision;
wire [17:0] value_variable_32_to_check;

wire enable_variable_32_to_check;
// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_32[5:0] = value_check_49_to_variable_32;
assign enable_check_to_variable_32[0] = enable_check_49_to_variable_32;
// 将变量节点32的输出与校验节点49的输入相连
assign value_variable_32_to_check_49 = value_variable_32_to_check[5:0];
assign enable_variable_32_to_check_49 = enable_variable_32_to_check;

// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_32[11:6] = value_check_50_to_variable_32;
assign enable_check_to_variable_32[1] = enable_check_50_to_variable_32;
// 将变量节点32的输出与校验节点50的输入相连
assign value_variable_32_to_check_50 = value_variable_32_to_check[11:6];
assign enable_variable_32_to_check_50 = enable_variable_32_to_check;

// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_32[17:12] = value_check_52_to_variable_32;
assign enable_check_to_variable_32[2] = enable_check_52_to_variable_32;
// 将变量节点32的输出与校验节点52的输入相连
assign value_variable_32_to_check_52 = value_variable_32_to_check[17:12];
assign enable_variable_32_to_check_52 = enable_variable_32_to_check;


// 变量节点33的接口
wire [17:0] value_check_to_variable_33;
wire [2:0] enable_check_to_variable_33;
wire [5:0] value_variable_33_to_decision;
wire [17:0] value_variable_33_to_check;

wire enable_variable_33_to_check;
// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_33[5:0] = value_check_53_to_variable_33;
assign enable_check_to_variable_33[0] = enable_check_53_to_variable_33;
// 将变量节点33的输出与校验节点53的输入相连
assign value_variable_33_to_check_53 = value_variable_33_to_check[5:0];
assign enable_variable_33_to_check_53 = enable_variable_33_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_33[11:6] = value_check_78_to_variable_33;
assign enable_check_to_variable_33[1] = enable_check_78_to_variable_33;
// 将变量节点33的输出与校验节点78的输入相连
assign value_variable_33_to_check_78 = value_variable_33_to_check[11:6];
assign enable_variable_33_to_check_78 = enable_variable_33_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_33[17:12] = value_check_122_to_variable_33;
assign enable_check_to_variable_33[2] = enable_check_122_to_variable_33;
// 将变量节点33的输出与校验节点122的输入相连
assign value_variable_33_to_check_122 = value_variable_33_to_check[17:12];
assign enable_variable_33_to_check_122 = enable_variable_33_to_check;


// 变量节点34的接口
wire [17:0] value_check_to_variable_34;
wire [2:0] enable_check_to_variable_34;
wire [5:0] value_variable_34_to_decision;
wire [17:0] value_variable_34_to_check;

wire enable_variable_34_to_check;
// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_34[5:0] = value_check_55_to_variable_34;
assign enable_check_to_variable_34[0] = enable_check_55_to_variable_34;
// 将变量节点34的输出与校验节点55的输入相连
assign value_variable_34_to_check_55 = value_variable_34_to_check[5:0];
assign enable_variable_34_to_check_55 = enable_variable_34_to_check;

// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_34[11:6] = value_check_98_to_variable_34;
assign enable_check_to_variable_34[1] = enable_check_98_to_variable_34;
// 将变量节点34的输出与校验节点98的输入相连
assign value_variable_34_to_check_98 = value_variable_34_to_check[11:6];
assign enable_variable_34_to_check_98 = enable_variable_34_to_check;

// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_34[17:12] = value_check_109_to_variable_34;
assign enable_check_to_variable_34[2] = enable_check_109_to_variable_34;
// 将变量节点34的输出与校验节点109的输入相连
assign value_variable_34_to_check_109 = value_variable_34_to_check[17:12];
assign enable_variable_34_to_check_109 = enable_variable_34_to_check;


// 变量节点35的接口
wire [17:0] value_check_to_variable_35;
wire [2:0] enable_check_to_variable_35;
wire [5:0] value_variable_35_to_decision;
wire [17:0] value_variable_35_to_check;

wire enable_variable_35_to_check;
// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_35[5:0] = value_check_58_to_variable_35;
assign enable_check_to_variable_35[0] = enable_check_58_to_variable_35;
// 将变量节点35的输出与校验节点58的输入相连
assign value_variable_35_to_check_58 = value_variable_35_to_check[5:0];
assign enable_variable_35_to_check_58 = enable_variable_35_to_check;

// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_35[11:6] = value_check_80_to_variable_35;
assign enable_check_to_variable_35[1] = enable_check_80_to_variable_35;
// 将变量节点35的输出与校验节点80的输入相连
assign value_variable_35_to_check_80 = value_variable_35_to_check[11:6];
assign enable_variable_35_to_check_80 = enable_variable_35_to_check;

// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_35[17:12] = value_check_86_to_variable_35;
assign enable_check_to_variable_35[2] = enable_check_86_to_variable_35;
// 将变量节点35的输出与校验节点86的输入相连
assign value_variable_35_to_check_86 = value_variable_35_to_check[17:12];
assign enable_variable_35_to_check_86 = enable_variable_35_to_check;


// 变量节点36的接口
wire [17:0] value_check_to_variable_36;
wire [2:0] enable_check_to_variable_36;
wire [5:0] value_variable_36_to_decision;
wire [17:0] value_variable_36_to_check;

wire enable_variable_36_to_check;
// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_36[5:0] = value_check_60_to_variable_36;
assign enable_check_to_variable_36[0] = enable_check_60_to_variable_36;
// 将变量节点36的输出与校验节点60的输入相连
assign value_variable_36_to_check_60 = value_variable_36_to_check[5:0];
assign enable_variable_36_to_check_60 = enable_variable_36_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_36[11:6] = value_check_112_to_variable_36;
assign enable_check_to_variable_36[1] = enable_check_112_to_variable_36;
// 将变量节点36的输出与校验节点112的输入相连
assign value_variable_36_to_check_112 = value_variable_36_to_check[11:6];
assign enable_variable_36_to_check_112 = enable_variable_36_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_36[17:12] = value_check_126_to_variable_36;
assign enable_check_to_variable_36[2] = enable_check_126_to_variable_36;
// 将变量节点36的输出与校验节点126的输入相连
assign value_variable_36_to_check_126 = value_variable_36_to_check[17:12];
assign enable_variable_36_to_check_126 = enable_variable_36_to_check;


// 变量节点37的接口
wire [17:0] value_check_to_variable_37;
wire [2:0] enable_check_to_variable_37;
wire [5:0] value_variable_37_to_decision;
wire [17:0] value_variable_37_to_check;

wire enable_variable_37_to_check;
// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_37[5:0] = value_check_64_to_variable_37;
assign enable_check_to_variable_37[0] = enable_check_64_to_variable_37;
// 将变量节点37的输出与校验节点64的输入相连
assign value_variable_37_to_check_64 = value_variable_37_to_check[5:0];
assign enable_variable_37_to_check_64 = enable_variable_37_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_37[11:6] = value_check_77_to_variable_37;
assign enable_check_to_variable_37[1] = enable_check_77_to_variable_37;
// 将变量节点37的输出与校验节点77的输入相连
assign value_variable_37_to_check_77 = value_variable_37_to_check[11:6];
assign enable_variable_37_to_check_77 = enable_variable_37_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_37[17:12] = value_check_89_to_variable_37;
assign enable_check_to_variable_37[2] = enable_check_89_to_variable_37;
// 将变量节点37的输出与校验节点89的输入相连
assign value_variable_37_to_check_89 = value_variable_37_to_check[17:12];
assign enable_variable_37_to_check_89 = enable_variable_37_to_check;


// 变量节点38的接口
wire [17:0] value_check_to_variable_38;
wire [2:0] enable_check_to_variable_38;
wire [5:0] value_variable_38_to_decision;
wire [17:0] value_variable_38_to_check;

wire enable_variable_38_to_check;
// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_38[5:0] = value_check_68_to_variable_38;
assign enable_check_to_variable_38[0] = enable_check_68_to_variable_38;
// 将变量节点38的输出与校验节点68的输入相连
assign value_variable_38_to_check_68 = value_variable_38_to_check[5:0];
assign enable_variable_38_to_check_68 = enable_variable_38_to_check;

// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_38[11:6] = value_check_69_to_variable_38;
assign enable_check_to_variable_38[1] = enable_check_69_to_variable_38;
// 将变量节点38的输出与校验节点69的输入相连
assign value_variable_38_to_check_69 = value_variable_38_to_check[11:6];
assign enable_variable_38_to_check_69 = enable_variable_38_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_38[17:12] = value_check_103_to_variable_38;
assign enable_check_to_variable_38[2] = enable_check_103_to_variable_38;
// 将变量节点38的输出与校验节点103的输入相连
assign value_variable_38_to_check_103 = value_variable_38_to_check[17:12];
assign enable_variable_38_to_check_103 = enable_variable_38_to_check;


// 变量节点39的接口
wire [17:0] value_check_to_variable_39;
wire [2:0] enable_check_to_variable_39;
wire [5:0] value_variable_39_to_decision;
wire [17:0] value_variable_39_to_check;

wire enable_variable_39_to_check;
// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_39[5:0] = value_check_70_to_variable_39;
assign enable_check_to_variable_39[0] = enable_check_70_to_variable_39;
// 将变量节点39的输出与校验节点70的输入相连
assign value_variable_39_to_check_70 = value_variable_39_to_check[5:0];
assign enable_variable_39_to_check_70 = enable_variable_39_to_check;

// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_39[11:6] = value_check_79_to_variable_39;
assign enable_check_to_variable_39[1] = enable_check_79_to_variable_39;
// 将变量节点39的输出与校验节点79的输入相连
assign value_variable_39_to_check_79 = value_variable_39_to_check[11:6];
assign enable_variable_39_to_check_79 = enable_variable_39_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_39[17:12] = value_check_118_to_variable_39;
assign enable_check_to_variable_39[2] = enable_check_118_to_variable_39;
// 将变量节点39的输出与校验节点118的输入相连
assign value_variable_39_to_check_118 = value_variable_39_to_check[17:12];
assign enable_variable_39_to_check_118 = enable_variable_39_to_check;


// 变量节点40的接口
wire [17:0] value_check_to_variable_40;
wire [2:0] enable_check_to_variable_40;
wire [5:0] value_variable_40_to_decision;
wire [17:0] value_variable_40_to_check;

wire enable_variable_40_to_check;
// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_40[5:0] = value_check_71_to_variable_40;
assign enable_check_to_variable_40[0] = enable_check_71_to_variable_40;
// 将变量节点40的输出与校验节点71的输入相连
assign value_variable_40_to_check_71 = value_variable_40_to_check[5:0];
assign enable_variable_40_to_check_71 = enable_variable_40_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_40[11:6] = value_check_92_to_variable_40;
assign enable_check_to_variable_40[1] = enable_check_92_to_variable_40;
// 将变量节点40的输出与校验节点92的输入相连
assign value_variable_40_to_check_92 = value_variable_40_to_check[11:6];
assign enable_variable_40_to_check_92 = enable_variable_40_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_40[17:12] = value_check_108_to_variable_40;
assign enable_check_to_variable_40[2] = enable_check_108_to_variable_40;
// 将变量节点40的输出与校验节点108的输入相连
assign value_variable_40_to_check_108 = value_variable_40_to_check[17:12];
assign enable_variable_40_to_check_108 = enable_variable_40_to_check;


// 变量节点41的接口
wire [17:0] value_check_to_variable_41;
wire [2:0] enable_check_to_variable_41;
wire [5:0] value_variable_41_to_decision;
wire [17:0] value_variable_41_to_check;

wire enable_variable_41_to_check;
// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_41[5:0] = value_check_82_to_variable_41;
assign enable_check_to_variable_41[0] = enable_check_82_to_variable_41;
// 将变量节点41的输出与校验节点82的输入相连
assign value_variable_41_to_check_82 = value_variable_41_to_check[5:0];
assign enable_variable_41_to_check_82 = enable_variable_41_to_check;

// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_41[11:6] = value_check_97_to_variable_41;
assign enable_check_to_variable_41[1] = enable_check_97_to_variable_41;
// 将变量节点41的输出与校验节点97的输入相连
assign value_variable_41_to_check_97 = value_variable_41_to_check[11:6];
assign enable_variable_41_to_check_97 = enable_variable_41_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_41[17:12] = value_check_102_to_variable_41;
assign enable_check_to_variable_41[2] = enable_check_102_to_variable_41;
// 将变量节点41的输出与校验节点102的输入相连
assign value_variable_41_to_check_102 = value_variable_41_to_check[17:12];
assign enable_variable_41_to_check_102 = enable_variable_41_to_check;


// 变量节点42的接口
wire [17:0] value_check_to_variable_42;
wire [2:0] enable_check_to_variable_42;
wire [5:0] value_variable_42_to_decision;
wire [17:0] value_variable_42_to_check;

wire enable_variable_42_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_42[5:0] = value_check_1_to_variable_42;
assign enable_check_to_variable_42[0] = enable_check_1_to_variable_42;
// 将变量节点42的输出与校验节点1的输入相连
assign value_variable_42_to_check_1 = value_variable_42_to_check[5:0];
assign enable_variable_42_to_check_1 = enable_variable_42_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_42[11:6] = value_check_115_to_variable_42;
assign enable_check_to_variable_42[1] = enable_check_115_to_variable_42;
// 将变量节点42的输出与校验节点115的输入相连
assign value_variable_42_to_check_115 = value_variable_42_to_check[11:6];
assign enable_variable_42_to_check_115 = enable_variable_42_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_42[17:12] = value_check_123_to_variable_42;
assign enable_check_to_variable_42[2] = enable_check_123_to_variable_42;
// 将变量节点42的输出与校验节点123的输入相连
assign value_variable_42_to_check_123 = value_variable_42_to_check[17:12];
assign enable_variable_42_to_check_123 = enable_variable_42_to_check;


// 变量节点43的接口
wire [17:0] value_check_to_variable_43;
wire [2:0] enable_check_to_variable_43;
wire [5:0] value_variable_43_to_decision;
wire [17:0] value_variable_43_to_check;

wire enable_variable_43_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_43[5:0] = value_check_0_to_variable_43;
assign enable_check_to_variable_43[0] = enable_check_0_to_variable_43;
// 将变量节点43的输出与校验节点0的输入相连
assign value_variable_43_to_check_0 = value_variable_43_to_check[5:0];
assign enable_variable_43_to_check_0 = enable_variable_43_to_check;

// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_43[11:6] = value_check_50_to_variable_43;
assign enable_check_to_variable_43[1] = enable_check_50_to_variable_43;
// 将变量节点43的输出与校验节点50的输入相连
assign value_variable_43_to_check_50 = value_variable_43_to_check[11:6];
assign enable_variable_43_to_check_50 = enable_variable_43_to_check;

// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_43[17:12] = value_check_80_to_variable_43;
assign enable_check_to_variable_43[2] = enable_check_80_to_variable_43;
// 将变量节点43的输出与校验节点80的输入相连
assign value_variable_43_to_check_80 = value_variable_43_to_check[17:12];
assign enable_variable_43_to_check_80 = enable_variable_43_to_check;


// 变量节点44的接口
wire [17:0] value_check_to_variable_44;
wire [2:0] enable_check_to_variable_44;
wire [5:0] value_variable_44_to_decision;
wire [17:0] value_variable_44_to_check;

wire enable_variable_44_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_44[5:0] = value_check_2_to_variable_44;
assign enable_check_to_variable_44[0] = enable_check_2_to_variable_44;
// 将变量节点44的输出与校验节点2的输入相连
assign value_variable_44_to_check_2 = value_variable_44_to_check[5:0];
assign enable_variable_44_to_check_2 = enable_variable_44_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_44[11:6] = value_check_61_to_variable_44;
assign enable_check_to_variable_44[1] = enable_check_61_to_variable_44;
// 将变量节点44的输出与校验节点61的输入相连
assign value_variable_44_to_check_61 = value_variable_44_to_check[11:6];
assign enable_variable_44_to_check_61 = enable_variable_44_to_check;

// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_44[17:12] = value_check_72_to_variable_44;
assign enable_check_to_variable_44[2] = enable_check_72_to_variable_44;
// 将变量节点44的输出与校验节点72的输入相连
assign value_variable_44_to_check_72 = value_variable_44_to_check[17:12];
assign enable_variable_44_to_check_72 = enable_variable_44_to_check;


// 变量节点45的接口
wire [17:0] value_check_to_variable_45;
wire [2:0] enable_check_to_variable_45;
wire [5:0] value_variable_45_to_decision;
wire [17:0] value_variable_45_to_check;

wire enable_variable_45_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_45[5:0] = value_check_3_to_variable_45;
assign enable_check_to_variable_45[0] = enable_check_3_to_variable_45;
// 将变量节点45的输出与校验节点3的输入相连
assign value_variable_45_to_check_3 = value_variable_45_to_check[5:0];
assign enable_variable_45_to_check_3 = enable_variable_45_to_check;

// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_45[11:6] = value_check_54_to_variable_45;
assign enable_check_to_variable_45[1] = enable_check_54_to_variable_45;
// 将变量节点45的输出与校验节点54的输入相连
assign value_variable_45_to_check_54 = value_variable_45_to_check[11:6];
assign enable_variable_45_to_check_54 = enable_variable_45_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_45[17:12] = value_check_96_to_variable_45;
assign enable_check_to_variable_45[2] = enable_check_96_to_variable_45;
// 将变量节点45的输出与校验节点96的输入相连
assign value_variable_45_to_check_96 = value_variable_45_to_check[17:12];
assign enable_variable_45_to_check_96 = enable_variable_45_to_check;


// 变量节点46的接口
wire [17:0] value_check_to_variable_46;
wire [2:0] enable_check_to_variable_46;
wire [5:0] value_variable_46_to_decision;
wire [17:0] value_variable_46_to_check;

wire enable_variable_46_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_46[5:0] = value_check_4_to_variable_46;
assign enable_check_to_variable_46[0] = enable_check_4_to_variable_46;
// 将变量节点46的输出与校验节点4的输入相连
assign value_variable_46_to_check_4 = value_variable_46_to_check[5:0];
assign enable_variable_46_to_check_4 = enable_variable_46_to_check;

// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_46[11:6] = value_check_20_to_variable_46;
assign enable_check_to_variable_46[1] = enable_check_20_to_variable_46;
// 将变量节点46的输出与校验节点20的输入相连
assign value_variable_46_to_check_20 = value_variable_46_to_check[11:6];
assign enable_variable_46_to_check_20 = enable_variable_46_to_check;

// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_46[17:12] = value_check_48_to_variable_46;
assign enable_check_to_variable_46[2] = enable_check_48_to_variable_46;
// 将变量节点46的输出与校验节点48的输入相连
assign value_variable_46_to_check_48 = value_variable_46_to_check[17:12];
assign enable_variable_46_to_check_48 = enable_variable_46_to_check;


// 变量节点47的接口
wire [17:0] value_check_to_variable_47;
wire [2:0] enable_check_to_variable_47;
wire [5:0] value_variable_47_to_decision;
wire [17:0] value_variable_47_to_check;

wire enable_variable_47_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_47[5:0] = value_check_5_to_variable_47;
assign enable_check_to_variable_47[0] = enable_check_5_to_variable_47;
// 将变量节点47的输出与校验节点5的输入相连
assign value_variable_47_to_check_5 = value_variable_47_to_check[5:0];
assign enable_variable_47_to_check_5 = enable_variable_47_to_check;

// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_47[11:6] = value_check_7_to_variable_47;
assign enable_check_to_variable_47[1] = enable_check_7_to_variable_47;
// 将变量节点47的输出与校验节点7的输入相连
assign value_variable_47_to_check_7 = value_variable_47_to_check[11:6];
assign enable_variable_47_to_check_7 = enable_variable_47_to_check;

// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_47[17:12] = value_check_86_to_variable_47;
assign enable_check_to_variable_47[2] = enable_check_86_to_variable_47;
// 将变量节点47的输出与校验节点86的输入相连
assign value_variable_47_to_check_86 = value_variable_47_to_check[17:12];
assign enable_variable_47_to_check_86 = enable_variable_47_to_check;


// 变量节点48的接口
wire [17:0] value_check_to_variable_48;
wire [2:0] enable_check_to_variable_48;
wire [5:0] value_variable_48_to_decision;
wire [17:0] value_variable_48_to_check;

wire enable_variable_48_to_check;
// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_48[5:0] = value_check_6_to_variable_48;
assign enable_check_to_variable_48[0] = enable_check_6_to_variable_48;
// 将变量节点48的输出与校验节点6的输入相连
assign value_variable_48_to_check_6 = value_variable_48_to_check[5:0];
assign enable_variable_48_to_check_6 = enable_variable_48_to_check;

// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_48[11:6] = value_check_69_to_variable_48;
assign enable_check_to_variable_48[1] = enable_check_69_to_variable_48;
// 将变量节点48的输出与校验节点69的输入相连
assign value_variable_48_to_check_69 = value_variable_48_to_check[11:6];
assign enable_variable_48_to_check_69 = enable_variable_48_to_check;

// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_48[17:12] = value_check_74_to_variable_48;
assign enable_check_to_variable_48[2] = enable_check_74_to_variable_48;
// 将变量节点48的输出与校验节点74的输入相连
assign value_variable_48_to_check_74 = value_variable_48_to_check[17:12];
assign enable_variable_48_to_check_74 = enable_variable_48_to_check;


// 变量节点49的接口
wire [17:0] value_check_to_variable_49;
wire [2:0] enable_check_to_variable_49;
wire [5:0] value_variable_49_to_decision;
wire [17:0] value_variable_49_to_check;

wire enable_variable_49_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_49[5:0] = value_check_8_to_variable_49;
assign enable_check_to_variable_49[0] = enable_check_8_to_variable_49;
// 将变量节点49的输出与校验节点8的输入相连
assign value_variable_49_to_check_8 = value_variable_49_to_check[5:0];
assign enable_variable_49_to_check_8 = enable_variable_49_to_check;

// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_49[11:6] = value_check_33_to_variable_49;
assign enable_check_to_variable_49[1] = enable_check_33_to_variable_49;
// 将变量节点49的输出与校验节点33的输入相连
assign value_variable_49_to_check_33 = value_variable_49_to_check[11:6];
assign enable_variable_49_to_check_33 = enable_variable_49_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_49[17:12] = value_check_78_to_variable_49;
assign enable_check_to_variable_49[2] = enable_check_78_to_variable_49;
// 将变量节点49的输出与校验节点78的输入相连
assign value_variable_49_to_check_78 = value_variable_49_to_check[17:12];
assign enable_variable_49_to_check_78 = enable_variable_49_to_check;


// 变量节点50的接口
wire [17:0] value_check_to_variable_50;
wire [2:0] enable_check_to_variable_50;
wire [5:0] value_variable_50_to_decision;
wire [17:0] value_variable_50_to_check;

wire enable_variable_50_to_check;
// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_50[5:0] = value_check_9_to_variable_50;
assign enable_check_to_variable_50[0] = enable_check_9_to_variable_50;
// 将变量节点50的输出与校验节点9的输入相连
assign value_variable_50_to_check_9 = value_variable_50_to_check[5:0];
assign enable_variable_50_to_check_9 = enable_variable_50_to_check;

// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_50[11:6] = value_check_25_to_variable_50;
assign enable_check_to_variable_50[1] = enable_check_25_to_variable_50;
// 将变量节点50的输出与校验节点25的输入相连
assign value_variable_50_to_check_25 = value_variable_50_to_check[11:6];
assign enable_variable_50_to_check_25 = enable_variable_50_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_50[17:12] = value_check_77_to_variable_50;
assign enable_check_to_variable_50[2] = enable_check_77_to_variable_50;
// 将变量节点50的输出与校验节点77的输入相连
assign value_variable_50_to_check_77 = value_variable_50_to_check[17:12];
assign enable_variable_50_to_check_77 = enable_variable_50_to_check;


// 变量节点51的接口
wire [17:0] value_check_to_variable_51;
wire [2:0] enable_check_to_variable_51;
wire [5:0] value_variable_51_to_decision;
wire [17:0] value_variable_51_to_check;

wire enable_variable_51_to_check;
// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_51[5:0] = value_check_10_to_variable_51;
assign enable_check_to_variable_51[0] = enable_check_10_to_variable_51;
// 将变量节点51的输出与校验节点10的输入相连
assign value_variable_51_to_check_10 = value_variable_51_to_check[5:0];
assign enable_variable_51_to_check_10 = enable_variable_51_to_check;

// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_51[11:6] = value_check_47_to_variable_51;
assign enable_check_to_variable_51[1] = enable_check_47_to_variable_51;
// 将变量节点51的输出与校验节点47的输入相连
assign value_variable_51_to_check_47 = value_variable_51_to_check[11:6];
assign enable_variable_51_to_check_47 = enable_variable_51_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_51[17:12] = value_check_122_to_variable_51;
assign enable_check_to_variable_51[2] = enable_check_122_to_variable_51;
// 将变量节点51的输出与校验节点122的输入相连
assign value_variable_51_to_check_122 = value_variable_51_to_check[17:12];
assign enable_variable_51_to_check_122 = enable_variable_51_to_check;


// 变量节点52的接口
wire [17:0] value_check_to_variable_52;
wire [2:0] enable_check_to_variable_52;
wire [5:0] value_variable_52_to_decision;
wire [17:0] value_variable_52_to_check;

wire enable_variable_52_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_52[5:0] = value_check_11_to_variable_52;
assign enable_check_to_variable_52[0] = enable_check_11_to_variable_52;
// 将变量节点52的输出与校验节点11的输入相连
assign value_variable_52_to_check_11 = value_variable_52_to_check[5:0];
assign enable_variable_52_to_check_11 = enable_variable_52_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_52[11:6] = value_check_34_to_variable_52;
assign enable_check_to_variable_52[1] = enable_check_34_to_variable_52;
// 将变量节点52的输出与校验节点34的输入相连
assign value_variable_52_to_check_34 = value_variable_52_to_check[11:6];
assign enable_variable_52_to_check_34 = enable_variable_52_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_52[17:12] = value_check_88_to_variable_52;
assign enable_check_to_variable_52[2] = enable_check_88_to_variable_52;
// 将变量节点52的输出与校验节点88的输入相连
assign value_variable_52_to_check_88 = value_variable_52_to_check[17:12];
assign enable_variable_52_to_check_88 = enable_variable_52_to_check;


// 变量节点53的接口
wire [17:0] value_check_to_variable_53;
wire [2:0] enable_check_to_variable_53;
wire [5:0] value_variable_53_to_decision;
wire [17:0] value_variable_53_to_check;

wire enable_variable_53_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_53[5:0] = value_check_12_to_variable_53;
assign enable_check_to_variable_53[0] = enable_check_12_to_variable_53;
// 将变量节点53的输出与校验节点12的输入相连
assign value_variable_53_to_check_12 = value_variable_53_to_check[5:0];
assign enable_variable_53_to_check_12 = enable_variable_53_to_check;

// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_53[11:6] = value_check_70_to_variable_53;
assign enable_check_to_variable_53[1] = enable_check_70_to_variable_53;
// 将变量节点53的输出与校验节点70的输入相连
assign value_variable_53_to_check_70 = value_variable_53_to_check[11:6];
assign enable_variable_53_to_check_70 = enable_variable_53_to_check;

// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_53[17:12] = value_check_110_to_variable_53;
assign enable_check_to_variable_53[2] = enable_check_110_to_variable_53;
// 将变量节点53的输出与校验节点110的输入相连
assign value_variable_53_to_check_110 = value_variable_53_to_check[17:12];
assign enable_variable_53_to_check_110 = enable_variable_53_to_check;


// 变量节点54的接口
wire [17:0] value_check_to_variable_54;
wire [2:0] enable_check_to_variable_54;
wire [5:0] value_variable_54_to_decision;
wire [17:0] value_variable_54_to_check;

wire enable_variable_54_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_54[5:0] = value_check_13_to_variable_54;
assign enable_check_to_variable_54[0] = enable_check_13_to_variable_54;
// 将变量节点54的输出与校验节点13的输入相连
assign value_variable_54_to_check_13 = value_variable_54_to_check[5:0];
assign enable_variable_54_to_check_13 = enable_variable_54_to_check;

// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_54[11:6] = value_check_97_to_variable_54;
assign enable_check_to_variable_54[1] = enable_check_97_to_variable_54;
// 将变量节点54的输出与校验节点97的输入相连
assign value_variable_54_to_check_97 = value_variable_54_to_check[11:6];
assign enable_variable_54_to_check_97 = enable_variable_54_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_54[17:12] = value_check_107_to_variable_54;
assign enable_check_to_variable_54[2] = enable_check_107_to_variable_54;
// 将变量节点54的输出与校验节点107的输入相连
assign value_variable_54_to_check_107 = value_variable_54_to_check[17:12];
assign enable_variable_54_to_check_107 = enable_variable_54_to_check;


// 变量节点55的接口
wire [17:0] value_check_to_variable_55;
wire [2:0] enable_check_to_variable_55;
wire [5:0] value_variable_55_to_decision;
wire [17:0] value_variable_55_to_check;

wire enable_variable_55_to_check;
// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_55[5:0] = value_check_14_to_variable_55;
assign enable_check_to_variable_55[0] = enable_check_14_to_variable_55;
// 将变量节点55的输出与校验节点14的输入相连
assign value_variable_55_to_check_14 = value_variable_55_to_check[5:0];
assign enable_variable_55_to_check_14 = enable_variable_55_to_check;

// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_55[11:6] = value_check_23_to_variable_55;
assign enable_check_to_variable_55[1] = enable_check_23_to_variable_55;
// 将变量节点55的输出与校验节点23的输入相连
assign value_variable_55_to_check_23 = value_variable_55_to_check[11:6];
assign enable_variable_55_to_check_23 = enable_variable_55_to_check;

// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_55[17:12] = value_check_83_to_variable_55;
assign enable_check_to_variable_55[2] = enable_check_83_to_variable_55;
// 将变量节点55的输出与校验节点83的输入相连
assign value_variable_55_to_check_83 = value_variable_55_to_check[17:12];
assign enable_variable_55_to_check_83 = enable_variable_55_to_check;


// 变量节点56的接口
wire [17:0] value_check_to_variable_56;
wire [2:0] enable_check_to_variable_56;
wire [5:0] value_variable_56_to_decision;
wire [17:0] value_variable_56_to_check;

wire enable_variable_56_to_check;
// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_56[5:0] = value_check_15_to_variable_56;
assign enable_check_to_variable_56[0] = enable_check_15_to_variable_56;
// 将变量节点56的输出与校验节点15的输入相连
assign value_variable_56_to_check_15 = value_variable_56_to_check[5:0];
assign enable_variable_56_to_check_15 = enable_variable_56_to_check;

// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_56[11:6] = value_check_46_to_variable_56;
assign enable_check_to_variable_56[1] = enable_check_46_to_variable_56;
// 将变量节点56的输出与校验节点46的输入相连
assign value_variable_56_to_check_46 = value_variable_56_to_check[11:6];
assign enable_variable_56_to_check_46 = enable_variable_56_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_56[17:12] = value_check_117_to_variable_56;
assign enable_check_to_variable_56[2] = enable_check_117_to_variable_56;
// 将变量节点56的输出与校验节点117的输入相连
assign value_variable_56_to_check_117 = value_variable_56_to_check[17:12];
assign enable_variable_56_to_check_117 = enable_variable_56_to_check;


// 变量节点57的接口
wire [17:0] value_check_to_variable_57;
wire [2:0] enable_check_to_variable_57;
wire [5:0] value_variable_57_to_decision;
wire [17:0] value_variable_57_to_check;

wire enable_variable_57_to_check;
// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_57[5:0] = value_check_16_to_variable_57;
assign enable_check_to_variable_57[0] = enable_check_16_to_variable_57;
// 将变量节点57的输出与校验节点16的输入相连
assign value_variable_57_to_check_16 = value_variable_57_to_check[5:0];
assign enable_variable_57_to_check_16 = enable_variable_57_to_check;

// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_57[11:6] = value_check_30_to_variable_57;
assign enable_check_to_variable_57[1] = enable_check_30_to_variable_57;
// 将变量节点57的输出与校验节点30的输入相连
assign value_variable_57_to_check_30 = value_variable_57_to_check[11:6];
assign enable_variable_57_to_check_30 = enable_variable_57_to_check;

// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_57[17:12] = value_check_62_to_variable_57;
assign enable_check_to_variable_57[2] = enable_check_62_to_variable_57;
// 将变量节点57的输出与校验节点62的输入相连
assign value_variable_57_to_check_62 = value_variable_57_to_check[17:12];
assign enable_variable_57_to_check_62 = enable_variable_57_to_check;


// 变量节点58的接口
wire [17:0] value_check_to_variable_58;
wire [2:0] enable_check_to_variable_58;
wire [5:0] value_variable_58_to_decision;
wire [17:0] value_variable_58_to_check;

wire enable_variable_58_to_check;
// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_58[5:0] = value_check_17_to_variable_58;
assign enable_check_to_variable_58[0] = enable_check_17_to_variable_58;
// 将变量节点58的输出与校验节点17的输入相连
assign value_variable_58_to_check_17 = value_variable_58_to_check[5:0];
assign enable_variable_58_to_check_17 = enable_variable_58_to_check;

// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_58[11:6] = value_check_52_to_variable_58;
assign enable_check_to_variable_58[1] = enable_check_52_to_variable_58;
// 将变量节点58的输出与校验节点52的输入相连
assign value_variable_58_to_check_52 = value_variable_58_to_check[11:6];
assign enable_variable_58_to_check_52 = enable_variable_58_to_check;

// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_58[17:12] = value_check_65_to_variable_58;
assign enable_check_to_variable_58[2] = enable_check_65_to_variable_58;
// 将变量节点58的输出与校验节点65的输入相连
assign value_variable_58_to_check_65 = value_variable_58_to_check[17:12];
assign enable_variable_58_to_check_65 = enable_variable_58_to_check;


// 变量节点59的接口
wire [17:0] value_check_to_variable_59;
wire [2:0] enable_check_to_variable_59;
wire [5:0] value_variable_59_to_decision;
wire [17:0] value_variable_59_to_check;

wire enable_variable_59_to_check;
// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_59[5:0] = value_check_18_to_variable_59;
assign enable_check_to_variable_59[0] = enable_check_18_to_variable_59;
// 将变量节点59的输出与校验节点18的输入相连
assign value_variable_59_to_check_18 = value_variable_59_to_check[5:0];
assign enable_variable_59_to_check_18 = enable_variable_59_to_check;

// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_59[11:6] = value_check_31_to_variable_59;
assign enable_check_to_variable_59[1] = enable_check_31_to_variable_59;
// 将变量节点59的输出与校验节点31的输入相连
assign value_variable_59_to_check_31 = value_variable_59_to_check[11:6];
assign enable_variable_59_to_check_31 = enable_variable_59_to_check;

// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_59[17:12] = value_check_95_to_variable_59;
assign enable_check_to_variable_59[2] = enable_check_95_to_variable_59;
// 将变量节点59的输出与校验节点95的输入相连
assign value_variable_59_to_check_95 = value_variable_59_to_check[17:12];
assign enable_variable_59_to_check_95 = enable_variable_59_to_check;


// 变量节点60的接口
wire [17:0] value_check_to_variable_60;
wire [2:0] enable_check_to_variable_60;
wire [5:0] value_variable_60_to_decision;
wire [17:0] value_variable_60_to_check;

wire enable_variable_60_to_check;
// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_60[5:0] = value_check_19_to_variable_60;
assign enable_check_to_variable_60[0] = enable_check_19_to_variable_60;
// 将变量节点60的输出与校验节点19的输入相连
assign value_variable_60_to_check_19 = value_variable_60_to_check[5:0];
assign enable_variable_60_to_check_19 = enable_variable_60_to_check;

// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_60[11:6] = value_check_56_to_variable_60;
assign enable_check_to_variable_60[1] = enable_check_56_to_variable_60;
// 将变量节点60的输出与校验节点56的输入相连
assign value_variable_60_to_check_56 = value_variable_60_to_check[11:6];
assign enable_variable_60_to_check_56 = enable_variable_60_to_check;

// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_60[17:12] = value_check_60_to_variable_60;
assign enable_check_to_variable_60[2] = enable_check_60_to_variable_60;
// 将变量节点60的输出与校验节点60的输入相连
assign value_variable_60_to_check_60 = value_variable_60_to_check[17:12];
assign enable_variable_60_to_check_60 = enable_variable_60_to_check;


// 变量节点61的接口
wire [17:0] value_check_to_variable_61;
wire [2:0] enable_check_to_variable_61;
wire [5:0] value_variable_61_to_decision;
wire [17:0] value_variable_61_to_check;

wire enable_variable_61_to_check;
// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_61[5:0] = value_check_21_to_variable_61;
assign enable_check_to_variable_61[0] = enable_check_21_to_variable_61;
// 将变量节点61的输出与校验节点21的输入相连
assign value_variable_61_to_check_21 = value_variable_61_to_check[5:0];
assign enable_variable_61_to_check_21 = enable_variable_61_to_check;

// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_61[11:6] = value_check_24_to_variable_61;
assign enable_check_to_variable_61[1] = enable_check_24_to_variable_61;
// 将变量节点61的输出与校验节点24的输入相连
assign value_variable_61_to_check_24 = value_variable_61_to_check[11:6];
assign enable_variable_61_to_check_24 = enable_variable_61_to_check;

// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_61[17:12] = value_check_71_to_variable_61;
assign enable_check_to_variable_61[2] = enable_check_71_to_variable_61;
// 将变量节点61的输出与校验节点71的输入相连
assign value_variable_61_to_check_71 = value_variable_61_to_check[17:12];
assign enable_variable_61_to_check_71 = enable_variable_61_to_check;


// 变量节点62的接口
wire [17:0] value_check_to_variable_62;
wire [2:0] enable_check_to_variable_62;
wire [5:0] value_variable_62_to_decision;
wire [17:0] value_variable_62_to_check;

wire enable_variable_62_to_check;
// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_62[5:0] = value_check_22_to_variable_62;
assign enable_check_to_variable_62[0] = enable_check_22_to_variable_62;
// 将变量节点62的输出与校验节点22的输入相连
assign value_variable_62_to_check_22 = value_variable_62_to_check[5:0];
assign enable_variable_62_to_check_22 = enable_variable_62_to_check;

// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_62[11:6] = value_check_45_to_variable_62;
assign enable_check_to_variable_62[1] = enable_check_45_to_variable_62;
// 将变量节点62的输出与校验节点45的输入相连
assign value_variable_62_to_check_45 = value_variable_62_to_check[11:6];
assign enable_variable_62_to_check_45 = enable_variable_62_to_check;

// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_62[17:12] = value_check_55_to_variable_62;
assign enable_check_to_variable_62[2] = enable_check_55_to_variable_62;
// 将变量节点62的输出与校验节点55的输入相连
assign value_variable_62_to_check_55 = value_variable_62_to_check[17:12];
assign enable_variable_62_to_check_55 = enable_variable_62_to_check;


// 变量节点63的接口
wire [17:0] value_check_to_variable_63;
wire [2:0] enable_check_to_variable_63;
wire [5:0] value_variable_63_to_decision;
wire [17:0] value_variable_63_to_check;

wire enable_variable_63_to_check;
// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_63[5:0] = value_check_26_to_variable_63;
assign enable_check_to_variable_63[0] = enable_check_26_to_variable_63;
// 将变量节点63的输出与校验节点26的输入相连
assign value_variable_63_to_check_26 = value_variable_63_to_check[5:0];
assign enable_variable_63_to_check_26 = enable_variable_63_to_check;

// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_63[11:6] = value_check_53_to_variable_63;
assign enable_check_to_variable_63[1] = enable_check_53_to_variable_63;
// 将变量节点63的输出与校验节点53的输入相连
assign value_variable_63_to_check_53 = value_variable_63_to_check[11:6];
assign enable_variable_63_to_check_53 = enable_variable_63_to_check;

// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_63[17:12] = value_check_76_to_variable_63;
assign enable_check_to_variable_63[2] = enable_check_76_to_variable_63;
// 将变量节点63的输出与校验节点76的输入相连
assign value_variable_63_to_check_76 = value_variable_63_to_check[17:12];
assign enable_variable_63_to_check_76 = enable_variable_63_to_check;


// 变量节点64的接口
wire [17:0] value_check_to_variable_64;
wire [2:0] enable_check_to_variable_64;
wire [5:0] value_variable_64_to_decision;
wire [17:0] value_variable_64_to_check;

wire enable_variable_64_to_check;
// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_64[5:0] = value_check_27_to_variable_64;
assign enable_check_to_variable_64[0] = enable_check_27_to_variable_64;
// 将变量节点64的输出与校验节点27的输入相连
assign value_variable_64_to_check_27 = value_variable_64_to_check[5:0];
assign enable_variable_64_to_check_27 = enable_variable_64_to_check;

// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_64[11:6] = value_check_35_to_variable_64;
assign enable_check_to_variable_64[1] = enable_check_35_to_variable_64;
// 将变量节点64的输出与校验节点35的输入相连
assign value_variable_64_to_check_35 = value_variable_64_to_check[11:6];
assign enable_variable_64_to_check_35 = enable_variable_64_to_check;

// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_64[17:12] = value_check_41_to_variable_64;
assign enable_check_to_variable_64[2] = enable_check_41_to_variable_64;
// 将变量节点64的输出与校验节点41的输入相连
assign value_variable_64_to_check_41 = value_variable_64_to_check[17:12];
assign enable_variable_64_to_check_41 = enable_variable_64_to_check;


// 变量节点65的接口
wire [17:0] value_check_to_variable_65;
wire [2:0] enable_check_to_variable_65;
wire [5:0] value_variable_65_to_decision;
wire [17:0] value_variable_65_to_check;

wire enable_variable_65_to_check;
// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_65[5:0] = value_check_28_to_variable_65;
assign enable_check_to_variable_65[0] = enable_check_28_to_variable_65;
// 将变量节点65的输出与校验节点28的输入相连
assign value_variable_65_to_check_28 = value_variable_65_to_check[5:0];
assign enable_variable_65_to_check_28 = enable_variable_65_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_65[11:6] = value_check_89_to_variable_65;
assign enable_check_to_variable_65[1] = enable_check_89_to_variable_65;
// 将变量节点65的输出与校验节点89的输入相连
assign value_variable_65_to_check_89 = value_variable_65_to_check[11:6];
assign enable_variable_65_to_check_89 = enable_variable_65_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_65[17:12] = value_check_124_to_variable_65;
assign enable_check_to_variable_65[2] = enable_check_124_to_variable_65;
// 将变量节点65的输出与校验节点124的输入相连
assign value_variable_65_to_check_124 = value_variable_65_to_check[17:12];
assign enable_variable_65_to_check_124 = enable_variable_65_to_check;


// 变量节点66的接口
wire [17:0] value_check_to_variable_66;
wire [2:0] enable_check_to_variable_66;
wire [5:0] value_variable_66_to_decision;
wire [17:0] value_variable_66_to_check;

wire enable_variable_66_to_check;
// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_66[5:0] = value_check_29_to_variable_66;
assign enable_check_to_variable_66[0] = enable_check_29_to_variable_66;
// 将变量节点66的输出与校验节点29的输入相连
assign value_variable_66_to_check_29 = value_variable_66_to_check[5:0];
assign enable_variable_66_to_check_29 = enable_variable_66_to_check;

// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_66[11:6] = value_check_44_to_variable_66;
assign enable_check_to_variable_66[1] = enable_check_44_to_variable_66;
// 将变量节点66的输出与校验节点44的输入相连
assign value_variable_66_to_check_44 = value_variable_66_to_check[11:6];
assign enable_variable_66_to_check_44 = enable_variable_66_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_66[17:12] = value_check_116_to_variable_66;
assign enable_check_to_variable_66[2] = enable_check_116_to_variable_66;
// 将变量节点66的输出与校验节点116的输入相连
assign value_variable_66_to_check_116 = value_variable_66_to_check[17:12];
assign enable_variable_66_to_check_116 = enable_variable_66_to_check;


// 变量节点67的接口
wire [17:0] value_check_to_variable_67;
wire [2:0] enable_check_to_variable_67;
wire [5:0] value_variable_67_to_decision;
wire [17:0] value_variable_67_to_check;

wire enable_variable_67_to_check;
// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_67[5:0] = value_check_32_to_variable_67;
assign enable_check_to_variable_67[0] = enable_check_32_to_variable_67;
// 将变量节点67的输出与校验节点32的输入相连
assign value_variable_67_to_check_32 = value_variable_67_to_check[5:0];
assign enable_variable_67_to_check_32 = enable_variable_67_to_check;

// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_67[11:6] = value_check_37_to_variable_67;
assign enable_check_to_variable_67[1] = enable_check_37_to_variable_67;
// 将变量节点67的输出与校验节点37的输入相连
assign value_variable_67_to_check_37 = value_variable_67_to_check[11:6];
assign enable_variable_67_to_check_37 = enable_variable_67_to_check;

// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_67[17:12] = value_check_98_to_variable_67;
assign enable_check_to_variable_67[2] = enable_check_98_to_variable_67;
// 将变量节点67的输出与校验节点98的输入相连
assign value_variable_67_to_check_98 = value_variable_67_to_check[17:12];
assign enable_variable_67_to_check_98 = enable_variable_67_to_check;


// 变量节点68的接口
wire [17:0] value_check_to_variable_68;
wire [2:0] enable_check_to_variable_68;
wire [5:0] value_variable_68_to_decision;
wire [17:0] value_variable_68_to_check;

wire enable_variable_68_to_check;
// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_68[5:0] = value_check_36_to_variable_68;
assign enable_check_to_variable_68[0] = enable_check_36_to_variable_68;
// 将变量节点68的输出与校验节点36的输入相连
assign value_variable_68_to_check_36 = value_variable_68_to_check[5:0];
assign enable_variable_68_to_check_36 = enable_variable_68_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_68[11:6] = value_check_84_to_variable_68;
assign enable_check_to_variable_68[1] = enable_check_84_to_variable_68;
// 将变量节点68的输出与校验节点84的输入相连
assign value_variable_68_to_check_84 = value_variable_68_to_check[11:6];
assign enable_variable_68_to_check_84 = enable_variable_68_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_68[17:12] = value_check_102_to_variable_68;
assign enable_check_to_variable_68[2] = enable_check_102_to_variable_68;
// 将变量节点68的输出与校验节点102的输入相连
assign value_variable_68_to_check_102 = value_variable_68_to_check[17:12];
assign enable_variable_68_to_check_102 = enable_variable_68_to_check;


// 变量节点69的接口
wire [17:0] value_check_to_variable_69;
wire [2:0] enable_check_to_variable_69;
wire [5:0] value_variable_69_to_decision;
wire [17:0] value_variable_69_to_check;

wire enable_variable_69_to_check;
// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_69[5:0] = value_check_38_to_variable_69;
assign enable_check_to_variable_69[0] = enable_check_38_to_variable_69;
// 将变量节点69的输出与校验节点38的输入相连
assign value_variable_69_to_check_38 = value_variable_69_to_check[5:0];
assign enable_variable_69_to_check_38 = enable_variable_69_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_69[11:6] = value_check_113_to_variable_69;
assign enable_check_to_variable_69[1] = enable_check_113_to_variable_69;
// 将变量节点69的输出与校验节点113的输入相连
assign value_variable_69_to_check_113 = value_variable_69_to_check[11:6];
assign enable_variable_69_to_check_113 = enable_variable_69_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_69[17:12] = value_check_115_to_variable_69;
assign enable_check_to_variable_69[2] = enable_check_115_to_variable_69;
// 将变量节点69的输出与校验节点115的输入相连
assign value_variable_69_to_check_115 = value_variable_69_to_check[17:12];
assign enable_variable_69_to_check_115 = enable_variable_69_to_check;


// 变量节点70的接口
wire [17:0] value_check_to_variable_70;
wire [2:0] enable_check_to_variable_70;
wire [5:0] value_variable_70_to_decision;
wire [17:0] value_variable_70_to_check;

wire enable_variable_70_to_check;
// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_70[5:0] = value_check_39_to_variable_70;
assign enable_check_to_variable_70[0] = enable_check_39_to_variable_70;
// 将变量节点70的输出与校验节点39的输入相连
assign value_variable_70_to_check_39 = value_variable_70_to_check[5:0];
assign enable_variable_70_to_check_39 = enable_variable_70_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_70[11:6] = value_check_92_to_variable_70;
assign enable_check_to_variable_70[1] = enable_check_92_to_variable_70;
// 将变量节点70的输出与校验节点92的输入相连
assign value_variable_70_to_check_92 = value_variable_70_to_check[11:6];
assign enable_variable_70_to_check_92 = enable_variable_70_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_70[17:12] = value_check_118_to_variable_70;
assign enable_check_to_variable_70[2] = enable_check_118_to_variable_70;
// 将变量节点70的输出与校验节点118的输入相连
assign value_variable_70_to_check_118 = value_variable_70_to_check[17:12];
assign enable_variable_70_to_check_118 = enable_variable_70_to_check;


// 变量节点71的接口
wire [17:0] value_check_to_variable_71;
wire [2:0] enable_check_to_variable_71;
wire [5:0] value_variable_71_to_decision;
wire [17:0] value_variable_71_to_check;

wire enable_variable_71_to_check;
// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_71[5:0] = value_check_40_to_variable_71;
assign enable_check_to_variable_71[0] = enable_check_40_to_variable_71;
// 将变量节点71的输出与校验节点40的输入相连
assign value_variable_71_to_check_40 = value_variable_71_to_check[5:0];
assign enable_variable_71_to_check_40 = enable_variable_71_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_71[11:6] = value_check_87_to_variable_71;
assign enable_check_to_variable_71[1] = enable_check_87_to_variable_71;
// 将变量节点71的输出与校验节点87的输入相连
assign value_variable_71_to_check_87 = value_variable_71_to_check[11:6];
assign enable_variable_71_to_check_87 = enable_variable_71_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_71[17:12] = value_check_91_to_variable_71;
assign enable_check_to_variable_71[2] = enable_check_91_to_variable_71;
// 将变量节点71的输出与校验节点91的输入相连
assign value_variable_71_to_check_91 = value_variable_71_to_check[17:12];
assign enable_variable_71_to_check_91 = enable_variable_71_to_check;


// 变量节点72的接口
wire [17:0] value_check_to_variable_72;
wire [2:0] enable_check_to_variable_72;
wire [5:0] value_variable_72_to_decision;
wire [17:0] value_variable_72_to_check;

wire enable_variable_72_to_check;
// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_72[5:0] = value_check_42_to_variable_72;
assign enable_check_to_variable_72[0] = enable_check_42_to_variable_72;
// 将变量节点72的输出与校验节点42的输入相连
assign value_variable_72_to_check_42 = value_variable_72_to_check[5:0];
assign enable_variable_72_to_check_42 = enable_variable_72_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_72[11:6] = value_check_93_to_variable_72;
assign enable_check_to_variable_72[1] = enable_check_93_to_variable_72;
// 将变量节点72的输出与校验节点93的输入相连
assign value_variable_72_to_check_93 = value_variable_72_to_check[11:6];
assign enable_variable_72_to_check_93 = enable_variable_72_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_72[17:12] = value_check_125_to_variable_72;
assign enable_check_to_variable_72[2] = enable_check_125_to_variable_72;
// 将变量节点72的输出与校验节点125的输入相连
assign value_variable_72_to_check_125 = value_variable_72_to_check[17:12];
assign enable_variable_72_to_check_125 = enable_variable_72_to_check;


// 变量节点73的接口
wire [17:0] value_check_to_variable_73;
wire [2:0] enable_check_to_variable_73;
wire [5:0] value_variable_73_to_decision;
wire [17:0] value_variable_73_to_check;

wire enable_variable_73_to_check;
// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_73[5:0] = value_check_43_to_variable_73;
assign enable_check_to_variable_73[0] = enable_check_43_to_variable_73;
// 将变量节点73的输出与校验节点43的输入相连
assign value_variable_73_to_check_43 = value_variable_73_to_check[5:0];
assign enable_variable_73_to_check_43 = enable_variable_73_to_check;

// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_73[11:6] = value_check_58_to_variable_73;
assign enable_check_to_variable_73[1] = enable_check_58_to_variable_73;
// 将变量节点73的输出与校验节点58的输入相连
assign value_variable_73_to_check_58 = value_variable_73_to_check[11:6];
assign enable_variable_73_to_check_58 = enable_variable_73_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_73[17:12] = value_check_103_to_variable_73;
assign enable_check_to_variable_73[2] = enable_check_103_to_variable_73;
// 将变量节点73的输出与校验节点103的输入相连
assign value_variable_73_to_check_103 = value_variable_73_to_check[17:12];
assign enable_variable_73_to_check_103 = enable_variable_73_to_check;


// 变量节点74的接口
wire [17:0] value_check_to_variable_74;
wire [2:0] enable_check_to_variable_74;
wire [5:0] value_variable_74_to_decision;
wire [17:0] value_variable_74_to_check;

wire enable_variable_74_to_check;
// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_74[5:0] = value_check_49_to_variable_74;
assign enable_check_to_variable_74[0] = enable_check_49_to_variable_74;
// 将变量节点74的输出与校验节点49的输入相连
assign value_variable_74_to_check_49 = value_variable_74_to_check[5:0];
assign enable_variable_74_to_check_49 = enable_variable_74_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_74[11:6] = value_check_111_to_variable_74;
assign enable_check_to_variable_74[1] = enable_check_111_to_variable_74;
// 将变量节点74的输出与校验节点111的输入相连
assign value_variable_74_to_check_111 = value_variable_74_to_check[11:6];
assign enable_variable_74_to_check_111 = enable_variable_74_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_74[17:12] = value_check_121_to_variable_74;
assign enable_check_to_variable_74[2] = enable_check_121_to_variable_74;
// 将变量节点74的输出与校验节点121的输入相连
assign value_variable_74_to_check_121 = value_variable_74_to_check[17:12];
assign enable_variable_74_to_check_121 = enable_variable_74_to_check;


// 变量节点75的接口
wire [17:0] value_check_to_variable_75;
wire [2:0] enable_check_to_variable_75;
wire [5:0] value_variable_75_to_decision;
wire [17:0] value_variable_75_to_check;

wire enable_variable_75_to_check;
// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_75[5:0] = value_check_51_to_variable_75;
assign enable_check_to_variable_75[0] = enable_check_51_to_variable_75;
// 将变量节点75的输出与校验节点51的输入相连
assign value_variable_75_to_check_51 = value_variable_75_to_check[5:0];
assign enable_variable_75_to_check_51 = enable_variable_75_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_75[11:6] = value_check_106_to_variable_75;
assign enable_check_to_variable_75[1] = enable_check_106_to_variable_75;
// 将变量节点75的输出与校验节点106的输入相连
assign value_variable_75_to_check_106 = value_variable_75_to_check[11:6];
assign enable_variable_75_to_check_106 = enable_variable_75_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_75[17:12] = value_check_120_to_variable_75;
assign enable_check_to_variable_75[2] = enable_check_120_to_variable_75;
// 将变量节点75的输出与校验节点120的输入相连
assign value_variable_75_to_check_120 = value_variable_75_to_check[17:12];
assign enable_variable_75_to_check_120 = enable_variable_75_to_check;


// 变量节点76的接口
wire [17:0] value_check_to_variable_76;
wire [2:0] enable_check_to_variable_76;
wire [5:0] value_variable_76_to_decision;
wire [17:0] value_variable_76_to_check;

wire enable_variable_76_to_check;
// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_76[5:0] = value_check_57_to_variable_76;
assign enable_check_to_variable_76[0] = enable_check_57_to_variable_76;
// 将变量节点76的输出与校验节点57的输入相连
assign value_variable_76_to_check_57 = value_variable_76_to_check[5:0];
assign enable_variable_76_to_check_57 = enable_variable_76_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_76[11:6] = value_check_81_to_variable_76;
assign enable_check_to_variable_76[1] = enable_check_81_to_variable_76;
// 将变量节点76的输出与校验节点81的输入相连
assign value_variable_76_to_check_81 = value_variable_76_to_check[11:6];
assign enable_variable_76_to_check_81 = enable_variable_76_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_76[17:12] = value_check_126_to_variable_76;
assign enable_check_to_variable_76[2] = enable_check_126_to_variable_76;
// 将变量节点76的输出与校验节点126的输入相连
assign value_variable_76_to_check_126 = value_variable_76_to_check[17:12];
assign enable_variable_76_to_check_126 = enable_variable_76_to_check;


// 变量节点77的接口
wire [17:0] value_check_to_variable_77;
wire [2:0] enable_check_to_variable_77;
wire [5:0] value_variable_77_to_decision;
wire [17:0] value_variable_77_to_check;

wire enable_variable_77_to_check;
// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_77[5:0] = value_check_59_to_variable_77;
assign enable_check_to_variable_77[0] = enable_check_59_to_variable_77;
// 将变量节点77的输出与校验节点59的输入相连
assign value_variable_77_to_check_59 = value_variable_77_to_check[5:0];
assign enable_variable_77_to_check_59 = enable_variable_77_to_check;

// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_77[11:6] = value_check_73_to_variable_77;
assign enable_check_to_variable_77[1] = enable_check_73_to_variable_77;
// 将变量节点77的输出与校验节点73的输入相连
assign value_variable_77_to_check_73 = value_variable_77_to_check[11:6];
assign enable_variable_77_to_check_73 = enable_variable_77_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_77[17:12] = value_check_85_to_variable_77;
assign enable_check_to_variable_77[2] = enable_check_85_to_variable_77;
// 将变量节点77的输出与校验节点85的输入相连
assign value_variable_77_to_check_85 = value_variable_77_to_check[17:12];
assign enable_variable_77_to_check_85 = enable_variable_77_to_check;


// 变量节点78的接口
wire [17:0] value_check_to_variable_78;
wire [2:0] enable_check_to_variable_78;
wire [5:0] value_variable_78_to_decision;
wire [17:0] value_variable_78_to_check;

wire enable_variable_78_to_check;
// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_78[5:0] = value_check_63_to_variable_78;
assign enable_check_to_variable_78[0] = enable_check_63_to_variable_78;
// 将变量节点78的输出与校验节点63的输入相连
assign value_variable_78_to_check_63 = value_variable_78_to_check[5:0];
assign enable_variable_78_to_check_63 = enable_variable_78_to_check;

// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_78[11:6] = value_check_68_to_variable_78;
assign enable_check_to_variable_78[1] = enable_check_68_to_variable_78;
// 将变量节点78的输出与校验节点68的输入相连
assign value_variable_78_to_check_68 = value_variable_78_to_check[11:6];
assign enable_variable_78_to_check_68 = enable_variable_78_to_check;

// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_78[17:12] = value_check_79_to_variable_78;
assign enable_check_to_variable_78[2] = enable_check_79_to_variable_78;
// 将变量节点78的输出与校验节点79的输入相连
assign value_variable_78_to_check_79 = value_variable_78_to_check[17:12];
assign enable_variable_78_to_check_79 = enable_variable_78_to_check;


// 变量节点79的接口
wire [17:0] value_check_to_variable_79;
wire [2:0] enable_check_to_variable_79;
wire [5:0] value_variable_79_to_decision;
wire [17:0] value_variable_79_to_check;

wire enable_variable_79_to_check;
// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_79[5:0] = value_check_64_to_variable_79;
assign enable_check_to_variable_79[0] = enable_check_64_to_variable_79;
// 将变量节点79的输出与校验节点64的输入相连
assign value_variable_79_to_check_64 = value_variable_79_to_check[5:0];
assign enable_variable_79_to_check_64 = enable_variable_79_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_79[11:6] = value_check_94_to_variable_79;
assign enable_check_to_variable_79[1] = enable_check_94_to_variable_79;
// 将变量节点79的输出与校验节点94的输入相连
assign value_variable_79_to_check_94 = value_variable_79_to_check[11:6];
assign enable_variable_79_to_check_94 = enable_variable_79_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_79[17:12] = value_check_119_to_variable_79;
assign enable_check_to_variable_79[2] = enable_check_119_to_variable_79;
// 将变量节点79的输出与校验节点119的输入相连
assign value_variable_79_to_check_119 = value_variable_79_to_check[17:12];
assign enable_variable_79_to_check_119 = enable_variable_79_to_check;


// 变量节点80的接口
wire [17:0] value_check_to_variable_80;
wire [2:0] enable_check_to_variable_80;
wire [5:0] value_variable_80_to_decision;
wire [17:0] value_variable_80_to_check;

wire enable_variable_80_to_check;
// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_80[5:0] = value_check_66_to_variable_80;
assign enable_check_to_variable_80[0] = enable_check_66_to_variable_80;
// 将变量节点80的输出与校验节点66的输入相连
assign value_variable_80_to_check_66 = value_variable_80_to_check[5:0];
assign enable_variable_80_to_check_66 = enable_variable_80_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_80[11:6] = value_check_101_to_variable_80;
assign enable_check_to_variable_80[1] = enable_check_101_to_variable_80;
// 将变量节点80的输出与校验节点101的输入相连
assign value_variable_80_to_check_101 = value_variable_80_to_check[11:6];
assign enable_variable_80_to_check_101 = enable_variable_80_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_80[17:12] = value_check_112_to_variable_80;
assign enable_check_to_variable_80[2] = enable_check_112_to_variable_80;
// 将变量节点80的输出与校验节点112的输入相连
assign value_variable_80_to_check_112 = value_variable_80_to_check[17:12];
assign enable_variable_80_to_check_112 = enable_variable_80_to_check;


// 变量节点81的接口
wire [17:0] value_check_to_variable_81;
wire [2:0] enable_check_to_variable_81;
wire [5:0] value_variable_81_to_decision;
wire [17:0] value_variable_81_to_check;

wire enable_variable_81_to_check;
// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_81[5:0] = value_check_67_to_variable_81;
assign enable_check_to_variable_81[0] = enable_check_67_to_variable_81;
// 将变量节点81的输出与校验节点67的输入相连
assign value_variable_81_to_check_67 = value_variable_81_to_check[5:0];
assign enable_variable_81_to_check_67 = enable_variable_81_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_81[11:6] = value_check_75_to_variable_81;
assign enable_check_to_variable_81[1] = enable_check_75_to_variable_81;
// 将变量节点81的输出与校验节点75的输入相连
assign value_variable_81_to_check_75 = value_variable_81_to_check[11:6];
assign enable_variable_81_to_check_75 = enable_variable_81_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_81[17:12] = value_check_108_to_variable_81;
assign enable_check_to_variable_81[2] = enable_check_108_to_variable_81;
// 将变量节点81的输出与校验节点108的输入相连
assign value_variable_81_to_check_108 = value_variable_81_to_check[17:12];
assign enable_variable_81_to_check_108 = enable_variable_81_to_check;


// 变量节点82的接口
wire [17:0] value_check_to_variable_82;
wire [2:0] enable_check_to_variable_82;
wire [5:0] value_variable_82_to_decision;
wire [17:0] value_variable_82_to_check;

wire enable_variable_82_to_check;
// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_82[5:0] = value_check_82_to_variable_82;
assign enable_check_to_variable_82[0] = enable_check_82_to_variable_82;
// 将变量节点82的输出与校验节点82的输入相连
assign value_variable_82_to_check_82 = value_variable_82_to_check[5:0];
assign enable_variable_82_to_check_82 = enable_variable_82_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_82[11:6] = value_check_90_to_variable_82;
assign enable_check_to_variable_82[1] = enable_check_90_to_variable_82;
// 将变量节点82的输出与校验节点90的输入相连
assign value_variable_82_to_check_90 = value_variable_82_to_check[11:6];
assign enable_variable_82_to_check_90 = enable_variable_82_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_82[17:12] = value_check_123_to_variable_82;
assign enable_check_to_variable_82[2] = enable_check_123_to_variable_82;
// 将变量节点82的输出与校验节点123的输入相连
assign value_variable_82_to_check_123 = value_variable_82_to_check[17:12];
assign enable_variable_82_to_check_123 = enable_variable_82_to_check;


// 变量节点83的接口
wire [17:0] value_check_to_variable_83;
wire [2:0] enable_check_to_variable_83;
wire [5:0] value_variable_83_to_decision;
wire [17:0] value_variable_83_to_check;

wire enable_variable_83_to_check;
// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_83[5:0] = value_check_99_to_variable_83;
assign enable_check_to_variable_83[0] = enable_check_99_to_variable_83;
// 将变量节点83的输出与校验节点99的输入相连
assign value_variable_83_to_check_99 = value_variable_83_to_check[5:0];
assign enable_variable_83_to_check_99 = enable_variable_83_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_83[11:6] = value_check_104_to_variable_83;
assign enable_check_to_variable_83[1] = enable_check_104_to_variable_83;
// 将变量节点83的输出与校验节点104的输入相连
assign value_variable_83_to_check_104 = value_variable_83_to_check[11:6];
assign enable_variable_83_to_check_104 = enable_variable_83_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_83[17:12] = value_check_105_to_variable_83;
assign enable_check_to_variable_83[2] = enable_check_105_to_variable_83;
// 将变量节点83的输出与校验节点105的输入相连
assign value_variable_83_to_check_105 = value_variable_83_to_check[17:12];
assign enable_variable_83_to_check_105 = enable_variable_83_to_check;


// 变量节点84的接口
wire [17:0] value_check_to_variable_84;
wire [2:0] enable_check_to_variable_84;
wire [5:0] value_variable_84_to_decision;
wire [17:0] value_variable_84_to_check;

wire enable_variable_84_to_check;
// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_84[5:0] = value_check_100_to_variable_84;
assign enable_check_to_variable_84[0] = enable_check_100_to_variable_84;
// 将变量节点84的输出与校验节点100的输入相连
assign value_variable_84_to_check_100 = value_variable_84_to_check[5:0];
assign enable_variable_84_to_check_100 = enable_variable_84_to_check;

// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_84[11:6] = value_check_110_to_variable_84;
assign enable_check_to_variable_84[1] = enable_check_110_to_variable_84;
// 将变量节点84的输出与校验节点110的输入相连
assign value_variable_84_to_check_110 = value_variable_84_to_check[11:6];
assign enable_variable_84_to_check_110 = enable_variable_84_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_84[17:12] = value_check_122_to_variable_84;
assign enable_check_to_variable_84[2] = enable_check_122_to_variable_84;
// 将变量节点84的输出与校验节点122的输入相连
assign value_variable_84_to_check_122 = value_variable_84_to_check[17:12];
assign enable_variable_84_to_check_122 = enable_variable_84_to_check;


// 变量节点85的接口
wire [17:0] value_check_to_variable_85;
wire [2:0] enable_check_to_variable_85;
wire [5:0] value_variable_85_to_decision;
wire [17:0] value_variable_85_to_check;

wire enable_variable_85_to_check;
// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_85[5:0] = value_check_109_to_variable_85;
assign enable_check_to_variable_85[0] = enable_check_109_to_variable_85;
// 将变量节点85的输出与校验节点109的输入相连
assign value_variable_85_to_check_109 = value_variable_85_to_check[5:0];
assign enable_variable_85_to_check_109 = enable_variable_85_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_85[11:6] = value_check_114_to_variable_85;
assign enable_check_to_variable_85[1] = enable_check_114_to_variable_85;
// 将变量节点85的输出与校验节点114的输入相连
assign value_variable_85_to_check_114 = value_variable_85_to_check[11:6];
assign enable_variable_85_to_check_114 = enable_variable_85_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_85[17:12] = value_check_127_to_variable_85;
assign enable_check_to_variable_85[2] = enable_check_127_to_variable_85;
// 将变量节点85的输出与校验节点127的输入相连
assign value_variable_85_to_check_127 = value_variable_85_to_check[17:12];
assign enable_variable_85_to_check_127 = enable_variable_85_to_check;


// 变量节点86的接口
wire [17:0] value_check_to_variable_86;
wire [2:0] enable_check_to_variable_86;
wire [5:0] value_variable_86_to_decision;
wire [17:0] value_variable_86_to_check;

wire enable_variable_86_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_86[5:0] = value_check_0_to_variable_86;
assign enable_check_to_variable_86[0] = enable_check_0_to_variable_86;
// 将变量节点86的输出与校验节点0的输入相连
assign value_variable_86_to_check_0 = value_variable_86_to_check[5:0];
assign enable_variable_86_to_check_0 = enable_variable_86_to_check;

// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_86[11:6] = value_check_57_to_variable_86;
assign enable_check_to_variable_86[1] = enable_check_57_to_variable_86;
// 将变量节点86的输出与校验节点57的输入相连
assign value_variable_86_to_check_57 = value_variable_86_to_check[11:6];
assign enable_variable_86_to_check_57 = enable_variable_86_to_check;

// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_86[17:12] = value_check_72_to_variable_86;
assign enable_check_to_variable_86[2] = enable_check_72_to_variable_86;
// 将变量节点86的输出与校验节点72的输入相连
assign value_variable_86_to_check_72 = value_variable_86_to_check[17:12];
assign enable_variable_86_to_check_72 = enable_variable_86_to_check;


// 变量节点87的接口
wire [17:0] value_check_to_variable_87;
wire [2:0] enable_check_to_variable_87;
wire [5:0] value_variable_87_to_decision;
wire [17:0] value_variable_87_to_check;

wire enable_variable_87_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_87[5:0] = value_check_1_to_variable_87;
assign enable_check_to_variable_87[0] = enable_check_1_to_variable_87;
// 将变量节点87的输出与校验节点1的输入相连
assign value_variable_87_to_check_1 = value_variable_87_to_check[5:0];
assign enable_variable_87_to_check_1 = enable_variable_87_to_check;

// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_87[11:6] = value_check_46_to_variable_87;
assign enable_check_to_variable_87[1] = enable_check_46_to_variable_87;
// 将变量节点87的输出与校验节点46的输入相连
assign value_variable_87_to_check_46 = value_variable_87_to_check[11:6];
assign enable_variable_87_to_check_46 = enable_variable_87_to_check;

// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_87[17:12] = value_check_48_to_variable_87;
assign enable_check_to_variable_87[2] = enable_check_48_to_variable_87;
// 将变量节点87的输出与校验节点48的输入相连
assign value_variable_87_to_check_48 = value_variable_87_to_check[17:12];
assign enable_variable_87_to_check_48 = enable_variable_87_to_check;


// 变量节点88的接口
wire [17:0] value_check_to_variable_88;
wire [2:0] enable_check_to_variable_88;
wire [5:0] value_variable_88_to_decision;
wire [17:0] value_variable_88_to_check;

wire enable_variable_88_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_88[5:0] = value_check_2_to_variable_88;
assign enable_check_to_variable_88[0] = enable_check_2_to_variable_88;
// 将变量节点88的输出与校验节点2的输入相连
assign value_variable_88_to_check_2 = value_variable_88_to_check[5:0];
assign enable_variable_88_to_check_2 = enable_variable_88_to_check;

// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_88[11:6] = value_check_68_to_variable_88;
assign enable_check_to_variable_88[1] = enable_check_68_to_variable_88;
// 将变量节点88的输出与校验节点68的输入相连
assign value_variable_88_to_check_68 = value_variable_88_to_check[11:6];
assign enable_variable_88_to_check_68 = enable_variable_88_to_check;

// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_88[17:12] = value_check_97_to_variable_88;
assign enable_check_to_variable_88[2] = enable_check_97_to_variable_88;
// 将变量节点88的输出与校验节点97的输入相连
assign value_variable_88_to_check_97 = value_variable_88_to_check[17:12];
assign enable_variable_88_to_check_97 = enable_variable_88_to_check;


// 变量节点89的接口
wire [17:0] value_check_to_variable_89;
wire [2:0] enable_check_to_variable_89;
wire [5:0] value_variable_89_to_decision;
wire [17:0] value_variable_89_to_check;

wire enable_variable_89_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_89[5:0] = value_check_3_to_variable_89;
assign enable_check_to_variable_89[0] = enable_check_3_to_variable_89;
// 将变量节点89的输出与校验节点3的输入相连
assign value_variable_89_to_check_3 = value_variable_89_to_check[5:0];
assign enable_variable_89_to_check_3 = enable_variable_89_to_check;

// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_89[11:6] = value_check_28_to_variable_89;
assign enable_check_to_variable_89[1] = enable_check_28_to_variable_89;
// 将变量节点89的输出与校验节点28的输入相连
assign value_variable_89_to_check_28 = value_variable_89_to_check[11:6];
assign enable_variable_89_to_check_28 = enable_variable_89_to_check;

// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_89[17:12] = value_check_36_to_variable_89;
assign enable_check_to_variable_89[2] = enable_check_36_to_variable_89;
// 将变量节点89的输出与校验节点36的输入相连
assign value_variable_89_to_check_36 = value_variable_89_to_check[17:12];
assign enable_variable_89_to_check_36 = enable_variable_89_to_check;


// 变量节点90的接口
wire [17:0] value_check_to_variable_90;
wire [2:0] enable_check_to_variable_90;
wire [5:0] value_variable_90_to_decision;
wire [17:0] value_variable_90_to_check;

wire enable_variable_90_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_90[5:0] = value_check_4_to_variable_90;
assign enable_check_to_variable_90[0] = enable_check_4_to_variable_90;
// 将变量节点90的输出与校验节点4的输入相连
assign value_variable_90_to_check_4 = value_variable_90_to_check[5:0];
assign enable_variable_90_to_check_4 = enable_variable_90_to_check;

// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_90[11:6] = value_check_41_to_variable_90;
assign enable_check_to_variable_90[1] = enable_check_41_to_variable_90;
// 将变量节点90的输出与校验节点41的输入相连
assign value_variable_90_to_check_41 = value_variable_90_to_check[11:6];
assign enable_variable_90_to_check_41 = enable_variable_90_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_90[17:12] = value_check_121_to_variable_90;
assign enable_check_to_variable_90[2] = enable_check_121_to_variable_90;
// 将变量节点90的输出与校验节点121的输入相连
assign value_variable_90_to_check_121 = value_variable_90_to_check[17:12];
assign enable_variable_90_to_check_121 = enable_variable_90_to_check;


// 变量节点91的接口
wire [17:0] value_check_to_variable_91;
wire [2:0] enable_check_to_variable_91;
wire [5:0] value_variable_91_to_decision;
wire [17:0] value_variable_91_to_check;

wire enable_variable_91_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_91[5:0] = value_check_5_to_variable_91;
assign enable_check_to_variable_91[0] = enable_check_5_to_variable_91;
// 将变量节点91的输出与校验节点5的输入相连
assign value_variable_91_to_check_5 = value_variable_91_to_check[5:0];
assign enable_variable_91_to_check_5 = enable_variable_91_to_check;

// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_91[11:6] = value_check_67_to_variable_91;
assign enable_check_to_variable_91[1] = enable_check_67_to_variable_91;
// 将变量节点91的输出与校验节点67的输入相连
assign value_variable_91_to_check_67 = value_variable_91_to_check[11:6];
assign enable_variable_91_to_check_67 = enable_variable_91_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_91[17:12] = value_check_112_to_variable_91;
assign enable_check_to_variable_91[2] = enable_check_112_to_variable_91;
// 将变量节点91的输出与校验节点112的输入相连
assign value_variable_91_to_check_112 = value_variable_91_to_check[17:12];
assign enable_variable_91_to_check_112 = enable_variable_91_to_check;


// 变量节点92的接口
wire [17:0] value_check_to_variable_92;
wire [2:0] enable_check_to_variable_92;
wire [5:0] value_variable_92_to_decision;
wire [17:0] value_variable_92_to_check;

wire enable_variable_92_to_check;
// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_92[5:0] = value_check_6_to_variable_92;
assign enable_check_to_variable_92[0] = enable_check_6_to_variable_92;
// 将变量节点92的输出与校验节点6的输入相连
assign value_variable_92_to_check_6 = value_variable_92_to_check[5:0];
assign enable_variable_92_to_check_6 = enable_variable_92_to_check;

// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_92[11:6] = value_check_19_to_variable_92;
assign enable_check_to_variable_92[1] = enable_check_19_to_variable_92;
// 将变量节点92的输出与校验节点19的输入相连
assign value_variable_92_to_check_19 = value_variable_92_to_check[11:6];
assign enable_variable_92_to_check_19 = enable_variable_92_to_check;

// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_92[17:12] = value_check_42_to_variable_92;
assign enable_check_to_variable_92[2] = enable_check_42_to_variable_92;
// 将变量节点92的输出与校验节点42的输入相连
assign value_variable_92_to_check_42 = value_variable_92_to_check[17:12];
assign enable_variable_92_to_check_42 = enable_variable_92_to_check;


// 变量节点93的接口
wire [17:0] value_check_to_variable_93;
wire [2:0] enable_check_to_variable_93;
wire [5:0] value_variable_93_to_decision;
wire [17:0] value_variable_93_to_check;

wire enable_variable_93_to_check;
// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_93[5:0] = value_check_7_to_variable_93;
assign enable_check_to_variable_93[0] = enable_check_7_to_variable_93;
// 将变量节点93的输出与校验节点7的输入相连
assign value_variable_93_to_check_7 = value_variable_93_to_check[5:0];
assign enable_variable_93_to_check_7 = enable_variable_93_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_93[11:6] = value_check_105_to_variable_93;
assign enable_check_to_variable_93[1] = enable_check_105_to_variable_93;
// 将变量节点93的输出与校验节点105的输入相连
assign value_variable_93_to_check_105 = value_variable_93_to_check[11:6];
assign enable_variable_93_to_check_105 = enable_variable_93_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_93[17:12] = value_check_118_to_variable_93;
assign enable_check_to_variable_93[2] = enable_check_118_to_variable_93;
// 将变量节点93的输出与校验节点118的输入相连
assign value_variable_93_to_check_118 = value_variable_93_to_check[17:12];
assign enable_variable_93_to_check_118 = enable_variable_93_to_check;


// 变量节点94的接口
wire [17:0] value_check_to_variable_94;
wire [2:0] enable_check_to_variable_94;
wire [5:0] value_variable_94_to_decision;
wire [17:0] value_variable_94_to_check;

wire enable_variable_94_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_94[5:0] = value_check_8_to_variable_94;
assign enable_check_to_variable_94[0] = enable_check_8_to_variable_94;
// 将变量节点94的输出与校验节点8的输入相连
assign value_variable_94_to_check_8 = value_variable_94_to_check[5:0];
assign enable_variable_94_to_check_8 = enable_variable_94_to_check;

// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_94[11:6] = value_check_23_to_variable_94;
assign enable_check_to_variable_94[1] = enable_check_23_to_variable_94;
// 将变量节点94的输出与校验节点23的输入相连
assign value_variable_94_to_check_23 = value_variable_94_to_check[11:6];
assign enable_variable_94_to_check_23 = enable_variable_94_to_check;

// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_94[17:12] = value_check_62_to_variable_94;
assign enable_check_to_variable_94[2] = enable_check_62_to_variable_94;
// 将变量节点94的输出与校验节点62的输入相连
assign value_variable_94_to_check_62 = value_variable_94_to_check[17:12];
assign enable_variable_94_to_check_62 = enable_variable_94_to_check;


// 变量节点95的接口
wire [17:0] value_check_to_variable_95;
wire [2:0] enable_check_to_variable_95;
wire [5:0] value_variable_95_to_decision;
wire [17:0] value_variable_95_to_check;

wire enable_variable_95_to_check;
// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_95[5:0] = value_check_9_to_variable_95;
assign enable_check_to_variable_95[0] = enable_check_9_to_variable_95;
// 将变量节点95的输出与校验节点9的输入相连
assign value_variable_95_to_check_9 = value_variable_95_to_check[5:0];
assign enable_variable_95_to_check_9 = enable_variable_95_to_check;

// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_95[11:6] = value_check_26_to_variable_95;
assign enable_check_to_variable_95[1] = enable_check_26_to_variable_95;
// 将变量节点95的输出与校验节点26的输入相连
assign value_variable_95_to_check_26 = value_variable_95_to_check[11:6];
assign enable_variable_95_to_check_26 = enable_variable_95_to_check;

// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_95[17:12] = value_check_98_to_variable_95;
assign enable_check_to_variable_95[2] = enable_check_98_to_variable_95;
// 将变量节点95的输出与校验节点98的输入相连
assign value_variable_95_to_check_98 = value_variable_95_to_check[17:12];
assign enable_variable_95_to_check_98 = enable_variable_95_to_check;


// 变量节点96的接口
wire [17:0] value_check_to_variable_96;
wire [2:0] enable_check_to_variable_96;
wire [5:0] value_variable_96_to_decision;
wire [17:0] value_variable_96_to_check;

wire enable_variable_96_to_check;
// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_96[5:0] = value_check_10_to_variable_96;
assign enable_check_to_variable_96[0] = enable_check_10_to_variable_96;
// 将变量节点96的输出与校验节点10的输入相连
assign value_variable_96_to_check_10 = value_variable_96_to_check[5:0];
assign enable_variable_96_to_check_10 = enable_variable_96_to_check;

// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_96[11:6] = value_check_22_to_variable_96;
assign enable_check_to_variable_96[1] = enable_check_22_to_variable_96;
// 将变量节点96的输出与校验节点22的输入相连
assign value_variable_96_to_check_22 = value_variable_96_to_check[11:6];
assign enable_variable_96_to_check_22 = enable_variable_96_to_check;

// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_96[17:12] = value_check_73_to_variable_96;
assign enable_check_to_variable_96[2] = enable_check_73_to_variable_96;
// 将变量节点96的输出与校验节点73的输入相连
assign value_variable_96_to_check_73 = value_variable_96_to_check[17:12];
assign enable_variable_96_to_check_73 = enable_variable_96_to_check;


// 变量节点97的接口
wire [17:0] value_check_to_variable_97;
wire [2:0] enable_check_to_variable_97;
wire [5:0] value_variable_97_to_decision;
wire [17:0] value_variable_97_to_check;

wire enable_variable_97_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_97[5:0] = value_check_11_to_variable_97;
assign enable_check_to_variable_97[0] = enable_check_11_to_variable_97;
// 将变量节点97的输出与校验节点11的输入相连
assign value_variable_97_to_check_11 = value_variable_97_to_check[5:0];
assign enable_variable_97_to_check_11 = enable_variable_97_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_97[11:6] = value_check_78_to_variable_97;
assign enable_check_to_variable_97[1] = enable_check_78_to_variable_97;
// 将变量节点97的输出与校验节点78的输入相连
assign value_variable_97_to_check_78 = value_variable_97_to_check[11:6];
assign enable_variable_97_to_check_78 = enable_variable_97_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_97[17:12] = value_check_126_to_variable_97;
assign enable_check_to_variable_97[2] = enable_check_126_to_variable_97;
// 将变量节点97的输出与校验节点126的输入相连
assign value_variable_97_to_check_126 = value_variable_97_to_check[17:12];
assign enable_variable_97_to_check_126 = enable_variable_97_to_check;


// 变量节点98的接口
wire [17:0] value_check_to_variable_98;
wire [2:0] enable_check_to_variable_98;
wire [5:0] value_variable_98_to_decision;
wire [17:0] value_variable_98_to_check;

wire enable_variable_98_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_98[5:0] = value_check_12_to_variable_98;
assign enable_check_to_variable_98[0] = enable_check_12_to_variable_98;
// 将变量节点98的输出与校验节点12的输入相连
assign value_variable_98_to_check_12 = value_variable_98_to_check[5:0];
assign enable_variable_98_to_check_12 = enable_variable_98_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_98[11:6] = value_check_87_to_variable_98;
assign enable_check_to_variable_98[1] = enable_check_87_to_variable_98;
// 将变量节点98的输出与校验节点87的输入相连
assign value_variable_98_to_check_87 = value_variable_98_to_check[11:6];
assign enable_variable_98_to_check_87 = enable_variable_98_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_98[17:12] = value_check_124_to_variable_98;
assign enable_check_to_variable_98[2] = enable_check_124_to_variable_98;
// 将变量节点98的输出与校验节点124的输入相连
assign value_variable_98_to_check_124 = value_variable_98_to_check[17:12];
assign enable_variable_98_to_check_124 = enable_variable_98_to_check;


// 变量节点99的接口
wire [17:0] value_check_to_variable_99;
wire [2:0] enable_check_to_variable_99;
wire [5:0] value_variable_99_to_decision;
wire [17:0] value_variable_99_to_check;

wire enable_variable_99_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_99[5:0] = value_check_13_to_variable_99;
assign enable_check_to_variable_99[0] = enable_check_13_to_variable_99;
// 将变量节点99的输出与校验节点13的输入相连
assign value_variable_99_to_check_13 = value_variable_99_to_check[5:0];
assign enable_variable_99_to_check_13 = enable_variable_99_to_check;

// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_99[11:6] = value_check_59_to_variable_99;
assign enable_check_to_variable_99[1] = enable_check_59_to_variable_99;
// 将变量节点99的输出与校验节点59的输入相连
assign value_variable_99_to_check_59 = value_variable_99_to_check[11:6];
assign enable_variable_99_to_check_59 = enable_variable_99_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_99[17:12] = value_check_101_to_variable_99;
assign enable_check_to_variable_99[2] = enable_check_101_to_variable_99;
// 将变量节点99的输出与校验节点101的输入相连
assign value_variable_99_to_check_101 = value_variable_99_to_check[17:12];
assign enable_variable_99_to_check_101 = enable_variable_99_to_check;


// 变量节点100的接口
wire [17:0] value_check_to_variable_100;
wire [2:0] enable_check_to_variable_100;
wire [5:0] value_variable_100_to_decision;
wire [17:0] value_variable_100_to_check;

wire enable_variable_100_to_check;
// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_100[5:0] = value_check_14_to_variable_100;
assign enable_check_to_variable_100[0] = enable_check_14_to_variable_100;
// 将变量节点100的输出与校验节点14的输入相连
assign value_variable_100_to_check_14 = value_variable_100_to_check[5:0];
assign enable_variable_100_to_check_14 = enable_variable_100_to_check;

// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_100[11:6] = value_check_57_to_variable_100;
assign enable_check_to_variable_100[1] = enable_check_57_to_variable_100;
// 将变量节点100的输出与校验节点57的输入相连
assign value_variable_100_to_check_57 = value_variable_100_to_check[11:6];
assign enable_variable_100_to_check_57 = enable_variable_100_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_100[17:12] = value_check_123_to_variable_100;
assign enable_check_to_variable_100[2] = enable_check_123_to_variable_100;
// 将变量节点100的输出与校验节点123的输入相连
assign value_variable_100_to_check_123 = value_variable_100_to_check[17:12];
assign enable_variable_100_to_check_123 = enable_variable_100_to_check;


// 变量节点101的接口
wire [17:0] value_check_to_variable_101;
wire [2:0] enable_check_to_variable_101;
wire [5:0] value_variable_101_to_decision;
wire [17:0] value_variable_101_to_check;

wire enable_variable_101_to_check;
// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_101[5:0] = value_check_15_to_variable_101;
assign enable_check_to_variable_101[0] = enable_check_15_to_variable_101;
// 将变量节点101的输出与校验节点15的输入相连
assign value_variable_101_to_check_15 = value_variable_101_to_check[5:0];
assign enable_variable_101_to_check_15 = enable_variable_101_to_check;

// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_101[11:6] = value_check_18_to_variable_101;
assign enable_check_to_variable_101[1] = enable_check_18_to_variable_101;
// 将变量节点101的输出与校验节点18的输入相连
assign value_variable_101_to_check_18 = value_variable_101_to_check[11:6];
assign enable_variable_101_to_check_18 = enable_variable_101_to_check;

// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_101[17:12] = value_check_37_to_variable_101;
assign enable_check_to_variable_101[2] = enable_check_37_to_variable_101;
// 将变量节点101的输出与校验节点37的输入相连
assign value_variable_101_to_check_37 = value_variable_101_to_check[17:12];
assign enable_variable_101_to_check_37 = enable_variable_101_to_check;


// 变量节点102的接口
wire [17:0] value_check_to_variable_102;
wire [2:0] enable_check_to_variable_102;
wire [5:0] value_variable_102_to_decision;
wire [17:0] value_variable_102_to_check;

wire enable_variable_102_to_check;
// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_102[5:0] = value_check_16_to_variable_102;
assign enable_check_to_variable_102[0] = enable_check_16_to_variable_102;
// 将变量节点102的输出与校验节点16的输入相连
assign value_variable_102_to_check_16 = value_variable_102_to_check[5:0];
assign enable_variable_102_to_check_16 = enable_variable_102_to_check;

// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_102[11:6] = value_check_17_to_variable_102;
assign enable_check_to_variable_102[1] = enable_check_17_to_variable_102;
// 将变量节点102的输出与校验节点17的输入相连
assign value_variable_102_to_check_17 = value_variable_102_to_check[11:6];
assign enable_variable_102_to_check_17 = enable_variable_102_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_102[17:12] = value_check_103_to_variable_102;
assign enable_check_to_variable_102[2] = enable_check_103_to_variable_102;
// 将变量节点102的输出与校验节点103的输入相连
assign value_variable_102_to_check_103 = value_variable_102_to_check[17:12];
assign enable_variable_102_to_check_103 = enable_variable_102_to_check;


// 变量节点103的接口
wire [17:0] value_check_to_variable_103;
wire [2:0] enable_check_to_variable_103;
wire [5:0] value_variable_103_to_decision;
wire [17:0] value_variable_103_to_check;

wire enable_variable_103_to_check;
// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_103[5:0] = value_check_20_to_variable_103;
assign enable_check_to_variable_103[0] = enable_check_20_to_variable_103;
// 将变量节点103的输出与校验节点20的输入相连
assign value_variable_103_to_check_20 = value_variable_103_to_check[5:0];
assign enable_variable_103_to_check_20 = enable_variable_103_to_check;

// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_103[11:6] = value_check_55_to_variable_103;
assign enable_check_to_variable_103[1] = enable_check_55_to_variable_103;
// 将变量节点103的输出与校验节点55的输入相连
assign value_variable_103_to_check_55 = value_variable_103_to_check[11:6];
assign enable_variable_103_to_check_55 = enable_variable_103_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_103[17:12] = value_check_75_to_variable_103;
assign enable_check_to_variable_103[2] = enable_check_75_to_variable_103;
// 将变量节点103的输出与校验节点75的输入相连
assign value_variable_103_to_check_75 = value_variable_103_to_check[17:12];
assign enable_variable_103_to_check_75 = enable_variable_103_to_check;


// 变量节点104的接口
wire [17:0] value_check_to_variable_104;
wire [2:0] enable_check_to_variable_104;
wire [5:0] value_variable_104_to_decision;
wire [17:0] value_variable_104_to_check;

wire enable_variable_104_to_check;
// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_104[5:0] = value_check_21_to_variable_104;
assign enable_check_to_variable_104[0] = enable_check_21_to_variable_104;
// 将变量节点104的输出与校验节点21的输入相连
assign value_variable_104_to_check_21 = value_variable_104_to_check[5:0];
assign enable_variable_104_to_check_21 = enable_variable_104_to_check;

// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_104[11:6] = value_check_29_to_variable_104;
assign enable_check_to_variable_104[1] = enable_check_29_to_variable_104;
// 将变量节点104的输出与校验节点29的输入相连
assign value_variable_104_to_check_29 = value_variable_104_to_check[11:6];
assign enable_variable_104_to_check_29 = enable_variable_104_to_check;

// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_104[17:12] = value_check_50_to_variable_104;
assign enable_check_to_variable_104[2] = enable_check_50_to_variable_104;
// 将变量节点104的输出与校验节点50的输入相连
assign value_variable_104_to_check_50 = value_variable_104_to_check[17:12];
assign enable_variable_104_to_check_50 = enable_variable_104_to_check;


// 变量节点105的接口
wire [17:0] value_check_to_variable_105;
wire [2:0] enable_check_to_variable_105;
wire [5:0] value_variable_105_to_decision;
wire [17:0] value_variable_105_to_check;

wire enable_variable_105_to_check;
// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_105[5:0] = value_check_24_to_variable_105;
assign enable_check_to_variable_105[0] = enable_check_24_to_variable_105;
// 将变量节点105的输出与校验节点24的输入相连
assign value_variable_105_to_check_24 = value_variable_105_to_check[5:0];
assign enable_variable_105_to_check_24 = enable_variable_105_to_check;

// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_105[11:6] = value_check_76_to_variable_105;
assign enable_check_to_variable_105[1] = enable_check_76_to_variable_105;
// 将变量节点105的输出与校验节点76的输入相连
assign value_variable_105_to_check_76 = value_variable_105_to_check[11:6];
assign enable_variable_105_to_check_76 = enable_variable_105_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_105[17:12] = value_check_119_to_variable_105;
assign enable_check_to_variable_105[2] = enable_check_119_to_variable_105;
// 将变量节点105的输出与校验节点119的输入相连
assign value_variable_105_to_check_119 = value_variable_105_to_check[17:12];
assign enable_variable_105_to_check_119 = enable_variable_105_to_check;


// 变量节点106的接口
wire [17:0] value_check_to_variable_106;
wire [2:0] enable_check_to_variable_106;
wire [5:0] value_variable_106_to_decision;
wire [17:0] value_variable_106_to_check;

wire enable_variable_106_to_check;
// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_106[5:0] = value_check_25_to_variable_106;
assign enable_check_to_variable_106[0] = enable_check_25_to_variable_106;
// 将变量节点106的输出与校验节点25的输入相连
assign value_variable_106_to_check_25 = value_variable_106_to_check[5:0];
assign enable_variable_106_to_check_25 = enable_variable_106_to_check;

// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_106[11:6] = value_check_44_to_variable_106;
assign enable_check_to_variable_106[1] = enable_check_44_to_variable_106;
// 将变量节点106的输出与校验节点44的输入相连
assign value_variable_106_to_check_44 = value_variable_106_to_check[11:6];
assign enable_variable_106_to_check_44 = enable_variable_106_to_check;

// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_106[17:12] = value_check_54_to_variable_106;
assign enable_check_to_variable_106[2] = enable_check_54_to_variable_106;
// 将变量节点106的输出与校验节点54的输入相连
assign value_variable_106_to_check_54 = value_variable_106_to_check[17:12];
assign enable_variable_106_to_check_54 = enable_variable_106_to_check;


// 变量节点107的接口
wire [17:0] value_check_to_variable_107;
wire [2:0] enable_check_to_variable_107;
wire [5:0] value_variable_107_to_decision;
wire [17:0] value_variable_107_to_check;

wire enable_variable_107_to_check;
// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_107[5:0] = value_check_27_to_variable_107;
assign enable_check_to_variable_107[0] = enable_check_27_to_variable_107;
// 将变量节点107的输出与校验节点27的输入相连
assign value_variable_107_to_check_27 = value_variable_107_to_check[5:0];
assign enable_variable_107_to_check_27 = enable_variable_107_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_107[11:6] = value_check_77_to_variable_107;
assign enable_check_to_variable_107[1] = enable_check_77_to_variable_107;
// 将变量节点107的输出与校验节点77的输入相连
assign value_variable_107_to_check_77 = value_variable_107_to_check[11:6];
assign enable_variable_107_to_check_77 = enable_variable_107_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_107[17:12] = value_check_113_to_variable_107;
assign enable_check_to_variable_107[2] = enable_check_113_to_variable_107;
// 将变量节点107的输出与校验节点113的输入相连
assign value_variable_107_to_check_113 = value_variable_107_to_check[17:12];
assign enable_variable_107_to_check_113 = enable_variable_107_to_check;


// 变量节点108的接口
wire [17:0] value_check_to_variable_108;
wire [2:0] enable_check_to_variable_108;
wire [5:0] value_variable_108_to_decision;
wire [17:0] value_variable_108_to_check;

wire enable_variable_108_to_check;
// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_108[5:0] = value_check_30_to_variable_108;
assign enable_check_to_variable_108[0] = enable_check_30_to_variable_108;
// 将变量节点108的输出与校验节点30的输入相连
assign value_variable_108_to_check_30 = value_variable_108_to_check[5:0];
assign enable_variable_108_to_check_30 = enable_variable_108_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_108[11:6] = value_check_92_to_variable_108;
assign enable_check_to_variable_108[1] = enable_check_92_to_variable_108;
// 将变量节点108的输出与校验节点92的输入相连
assign value_variable_108_to_check_92 = value_variable_108_to_check[11:6];
assign enable_variable_108_to_check_92 = enable_variable_108_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_108[17:12] = value_check_111_to_variable_108;
assign enable_check_to_variable_108[2] = enable_check_111_to_variable_108;
// 将变量节点108的输出与校验节点111的输入相连
assign value_variable_108_to_check_111 = value_variable_108_to_check[17:12];
assign enable_variable_108_to_check_111 = enable_variable_108_to_check;


// 变量节点109的接口
wire [17:0] value_check_to_variable_109;
wire [2:0] enable_check_to_variable_109;
wire [5:0] value_variable_109_to_decision;
wire [17:0] value_variable_109_to_check;

wire enable_variable_109_to_check;
// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_109[5:0] = value_check_31_to_variable_109;
assign enable_check_to_variable_109[0] = enable_check_31_to_variable_109;
// 将变量节点109的输出与校验节点31的输入相连
assign value_variable_109_to_check_31 = value_variable_109_to_check[5:0];
assign enable_variable_109_to_check_31 = enable_variable_109_to_check;

// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_109[11:6] = value_check_58_to_variable_109;
assign enable_check_to_variable_109[1] = enable_check_58_to_variable_109;
// 将变量节点109的输出与校验节点58的输入相连
assign value_variable_109_to_check_58 = value_variable_109_to_check[11:6];
assign enable_variable_109_to_check_58 = enable_variable_109_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_109[17:12] = value_check_78_to_variable_109;
assign enable_check_to_variable_109[2] = enable_check_78_to_variable_109;
// 将变量节点109的输出与校验节点78的输入相连
assign value_variable_109_to_check_78 = value_variable_109_to_check[17:12];
assign enable_variable_109_to_check_78 = enable_variable_109_to_check;


// 变量节点110的接口
wire [17:0] value_check_to_variable_110;
wire [2:0] enable_check_to_variable_110;
wire [5:0] value_variable_110_to_decision;
wire [17:0] value_variable_110_to_check;

wire enable_variable_110_to_check;
// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_110[5:0] = value_check_32_to_variable_110;
assign enable_check_to_variable_110[0] = enable_check_32_to_variable_110;
// 将变量节点110的输出与校验节点32的输入相连
assign value_variable_110_to_check_32 = value_variable_110_to_check[5:0];
assign enable_variable_110_to_check_32 = enable_variable_110_to_check;

// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_110[11:6] = value_check_69_to_variable_110;
assign enable_check_to_variable_110[1] = enable_check_69_to_variable_110;
// 将变量节点110的输出与校验节点69的输入相连
assign value_variable_110_to_check_69 = value_variable_110_to_check[11:6];
assign enable_variable_110_to_check_69 = enable_variable_110_to_check;

// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_110[17:12] = value_check_71_to_variable_110;
assign enable_check_to_variable_110[2] = enable_check_71_to_variable_110;
// 将变量节点110的输出与校验节点71的输入相连
assign value_variable_110_to_check_71 = value_variable_110_to_check[17:12];
assign enable_variable_110_to_check_71 = enable_variable_110_to_check;


// 变量节点111的接口
wire [17:0] value_check_to_variable_111;
wire [2:0] enable_check_to_variable_111;
wire [5:0] value_variable_111_to_decision;
wire [17:0] value_variable_111_to_check;

wire enable_variable_111_to_check;
// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_111[5:0] = value_check_33_to_variable_111;
assign enable_check_to_variable_111[0] = enable_check_33_to_variable_111;
// 将变量节点111的输出与校验节点33的输入相连
assign value_variable_111_to_check_33 = value_variable_111_to_check[5:0];
assign enable_variable_111_to_check_33 = enable_variable_111_to_check;

// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_111[11:6] = value_check_64_to_variable_111;
assign enable_check_to_variable_111[1] = enable_check_64_to_variable_111;
// 将变量节点111的输出与校验节点64的输入相连
assign value_variable_111_to_check_64 = value_variable_111_to_check[11:6];
assign enable_variable_111_to_check_64 = enable_variable_111_to_check;

// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_111[17:12] = value_check_79_to_variable_111;
assign enable_check_to_variable_111[2] = enable_check_79_to_variable_111;
// 将变量节点111的输出与校验节点79的输入相连
assign value_variable_111_to_check_79 = value_variable_111_to_check[17:12];
assign enable_variable_111_to_check_79 = enable_variable_111_to_check;


// 变量节点112的接口
wire [17:0] value_check_to_variable_112;
wire [2:0] enable_check_to_variable_112;
wire [5:0] value_variable_112_to_decision;
wire [17:0] value_variable_112_to_check;

wire enable_variable_112_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_112[5:0] = value_check_12_to_variable_112;
assign enable_check_to_variable_112[0] = enable_check_12_to_variable_112;
// 将变量节点112的输出与校验节点12的输入相连
assign value_variable_112_to_check_12 = value_variable_112_to_check[5:0];
assign enable_variable_112_to_check_12 = enable_variable_112_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_112[11:6] = value_check_34_to_variable_112;
assign enable_check_to_variable_112[1] = enable_check_34_to_variable_112;
// 将变量节点112的输出与校验节点34的输入相连
assign value_variable_112_to_check_34 = value_variable_112_to_check[11:6];
assign enable_variable_112_to_check_34 = enable_variable_112_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_112[17:12] = value_check_90_to_variable_112;
assign enable_check_to_variable_112[2] = enable_check_90_to_variable_112;
// 将变量节点112的输出与校验节点90的输入相连
assign value_variable_112_to_check_90 = value_variable_112_to_check[17:12];
assign enable_variable_112_to_check_90 = enable_variable_112_to_check;


// 变量节点113的接口
wire [17:0] value_check_to_variable_113;
wire [2:0] enable_check_to_variable_113;
wire [5:0] value_variable_113_to_decision;
wire [17:0] value_variable_113_to_check;

wire enable_variable_113_to_check;
// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_113[5:0] = value_check_35_to_variable_113;
assign enable_check_to_variable_113[0] = enable_check_35_to_variable_113;
// 将变量节点113的输出与校验节点35的输入相连
assign value_variable_113_to_check_35 = value_variable_113_to_check[5:0];
assign enable_variable_113_to_check_35 = enable_variable_113_to_check;

// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_113[11:6] = value_check_63_to_variable_113;
assign enable_check_to_variable_113[1] = enable_check_63_to_variable_113;
// 将变量节点113的输出与校验节点63的输入相连
assign value_variable_113_to_check_63 = value_variable_113_to_check[11:6];
assign enable_variable_113_to_check_63 = enable_variable_113_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_113[17:12] = value_check_120_to_variable_113;
assign enable_check_to_variable_113[2] = enable_check_120_to_variable_113;
// 将变量节点113的输出与校验节点120的输入相连
assign value_variable_113_to_check_120 = value_variable_113_to_check[17:12];
assign enable_variable_113_to_check_120 = enable_variable_113_to_check;


// 变量节点114的接口
wire [17:0] value_check_to_variable_114;
wire [2:0] enable_check_to_variable_114;
wire [5:0] value_variable_114_to_decision;
wire [17:0] value_variable_114_to_check;

wire enable_variable_114_to_check;
// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_114[5:0] = value_check_38_to_variable_114;
assign enable_check_to_variable_114[0] = enable_check_38_to_variable_114;
// 将变量节点114的输出与校验节点38的输入相连
assign value_variable_114_to_check_38 = value_variable_114_to_check[5:0];
assign enable_variable_114_to_check_38 = enable_variable_114_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_114[11:6] = value_check_61_to_variable_114;
assign enable_check_to_variable_114[1] = enable_check_61_to_variable_114;
// 将变量节点114的输出与校验节点61的输入相连
assign value_variable_114_to_check_61 = value_variable_114_to_check[11:6];
assign enable_variable_114_to_check_61 = enable_variable_114_to_check;

// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_114[17:12] = value_check_65_to_variable_114;
assign enable_check_to_variable_114[2] = enable_check_65_to_variable_114;
// 将变量节点114的输出与校验节点65的输入相连
assign value_variable_114_to_check_65 = value_variable_114_to_check[17:12];
assign enable_variable_114_to_check_65 = enable_variable_114_to_check;


// 变量节点115的接口
wire [17:0] value_check_to_variable_115;
wire [2:0] enable_check_to_variable_115;
wire [5:0] value_variable_115_to_decision;
wire [17:0] value_variable_115_to_check;

wire enable_variable_115_to_check;
// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_115[5:0] = value_check_39_to_variable_115;
assign enable_check_to_variable_115[0] = enable_check_39_to_variable_115;
// 将变量节点115的输出与校验节点39的输入相连
assign value_variable_115_to_check_39 = value_variable_115_to_check[5:0];
assign enable_variable_115_to_check_39 = enable_variable_115_to_check;

// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_115[11:6] = value_check_100_to_variable_115;
assign enable_check_to_variable_115[1] = enable_check_100_to_variable_115;
// 将变量节点115的输出与校验节点100的输入相连
assign value_variable_115_to_check_100 = value_variable_115_to_check[11:6];
assign enable_variable_115_to_check_100 = enable_variable_115_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_115[17:12] = value_check_102_to_variable_115;
assign enable_check_to_variable_115[2] = enable_check_102_to_variable_115;
// 将变量节点115的输出与校验节点102的输入相连
assign value_variable_115_to_check_102 = value_variable_115_to_check[17:12];
assign enable_variable_115_to_check_102 = enable_variable_115_to_check;


// 变量节点116的接口
wire [17:0] value_check_to_variable_116;
wire [2:0] enable_check_to_variable_116;
wire [5:0] value_variable_116_to_decision;
wire [17:0] value_variable_116_to_check;

wire enable_variable_116_to_check;
// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_116[5:0] = value_check_40_to_variable_116;
assign enable_check_to_variable_116[0] = enable_check_40_to_variable_116;
// 将变量节点116的输出与校验节点40的输入相连
assign value_variable_116_to_check_40 = value_variable_116_to_check[5:0];
assign enable_variable_116_to_check_40 = enable_variable_116_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_116[11:6] = value_check_84_to_variable_116;
assign enable_check_to_variable_116[1] = enable_check_84_to_variable_116;
// 将变量节点116的输出与校验节点84的输入相连
assign value_variable_116_to_check_84 = value_variable_116_to_check[11:6];
assign enable_variable_116_to_check_84 = enable_variable_116_to_check;

// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_116[17:12] = value_check_109_to_variable_116;
assign enable_check_to_variable_116[2] = enable_check_109_to_variable_116;
// 将变量节点116的输出与校验节点109的输入相连
assign value_variable_116_to_check_109 = value_variable_116_to_check[17:12];
assign enable_variable_116_to_check_109 = enable_variable_116_to_check;


// 变量节点117的接口
wire [17:0] value_check_to_variable_117;
wire [2:0] enable_check_to_variable_117;
wire [5:0] value_variable_117_to_decision;
wire [17:0] value_variable_117_to_check;

wire enable_variable_117_to_check;
// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_117[5:0] = value_check_43_to_variable_117;
assign enable_check_to_variable_117[0] = enable_check_43_to_variable_117;
// 将变量节点117的输出与校验节点43的输入相连
assign value_variable_117_to_check_43 = value_variable_117_to_check[5:0];
assign enable_variable_117_to_check_43 = enable_variable_117_to_check;

// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_117[11:6] = value_check_56_to_variable_117;
assign enable_check_to_variable_117[1] = enable_check_56_to_variable_117;
// 将变量节点117的输出与校验节点56的输入相连
assign value_variable_117_to_check_56 = value_variable_117_to_check[11:6];
assign enable_variable_117_to_check_56 = enable_variable_117_to_check;

// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_117[17:12] = value_check_99_to_variable_117;
assign enable_check_to_variable_117[2] = enable_check_99_to_variable_117;
// 将变量节点117的输出与校验节点99的输入相连
assign value_variable_117_to_check_99 = value_variable_117_to_check[17:12];
assign enable_variable_117_to_check_99 = enable_variable_117_to_check;


// 变量节点118的接口
wire [17:0] value_check_to_variable_118;
wire [2:0] enable_check_to_variable_118;
wire [5:0] value_variable_118_to_decision;
wire [17:0] value_variable_118_to_check;

wire enable_variable_118_to_check;
// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_118[5:0] = value_check_45_to_variable_118;
assign enable_check_to_variable_118[0] = enable_check_45_to_variable_118;
// 将变量节点118的输出与校验节点45的输入相连
assign value_variable_118_to_check_45 = value_variable_118_to_check[5:0];
assign enable_variable_118_to_check_45 = enable_variable_118_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_118[11:6] = value_check_93_to_variable_118;
assign enable_check_to_variable_118[1] = enable_check_93_to_variable_118;
// 将变量节点118的输出与校验节点93的输入相连
assign value_variable_118_to_check_93 = value_variable_118_to_check[11:6];
assign enable_variable_118_to_check_93 = enable_variable_118_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_118[17:12] = value_check_107_to_variable_118;
assign enable_check_to_variable_118[2] = enable_check_107_to_variable_118;
// 将变量节点118的输出与校验节点107的输入相连
assign value_variable_118_to_check_107 = value_variable_118_to_check[17:12];
assign enable_variable_118_to_check_107 = enable_variable_118_to_check;


// 变量节点119的接口
wire [17:0] value_check_to_variable_119;
wire [2:0] enable_check_to_variable_119;
wire [5:0] value_variable_119_to_decision;
wire [17:0] value_variable_119_to_check;

wire enable_variable_119_to_check;
// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_119[5:0] = value_check_47_to_variable_119;
assign enable_check_to_variable_119[0] = enable_check_47_to_variable_119;
// 将变量节点119的输出与校验节点47的输入相连
assign value_variable_119_to_check_47 = value_variable_119_to_check[5:0];
assign enable_variable_119_to_check_47 = enable_variable_119_to_check;

// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_119[11:6] = value_check_49_to_variable_119;
assign enable_check_to_variable_119[1] = enable_check_49_to_variable_119;
// 将变量节点119的输出与校验节点49的输入相连
assign value_variable_119_to_check_49 = value_variable_119_to_check[11:6];
assign enable_variable_119_to_check_49 = enable_variable_119_to_check;

// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_119[17:12] = value_check_51_to_variable_119;
assign enable_check_to_variable_119[2] = enable_check_51_to_variable_119;
// 将变量节点119的输出与校验节点51的输入相连
assign value_variable_119_to_check_51 = value_variable_119_to_check[17:12];
assign enable_variable_119_to_check_51 = enable_variable_119_to_check;


// 变量节点120的接口
wire [17:0] value_check_to_variable_120;
wire [2:0] enable_check_to_variable_120;
wire [5:0] value_variable_120_to_decision;
wire [17:0] value_variable_120_to_check;

wire enable_variable_120_to_check;
// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_120[5:0] = value_check_52_to_variable_120;
assign enable_check_to_variable_120[0] = enable_check_52_to_variable_120;
// 将变量节点120的输出与校验节点52的输入相连
assign value_variable_120_to_check_52 = value_variable_120_to_check[5:0];
assign enable_variable_120_to_check_52 = enable_variable_120_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_120[11:6] = value_check_94_to_variable_120;
assign enable_check_to_variable_120[1] = enable_check_94_to_variable_120;
// 将变量节点120的输出与校验节点94的输入相连
assign value_variable_120_to_check_94 = value_variable_120_to_check[11:6];
assign enable_variable_120_to_check_94 = enable_variable_120_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_120[17:12] = value_check_114_to_variable_120;
assign enable_check_to_variable_120[2] = enable_check_114_to_variable_120;
// 将变量节点120的输出与校验节点114的输入相连
assign value_variable_120_to_check_114 = value_variable_120_to_check[17:12];
assign enable_variable_120_to_check_114 = enable_variable_120_to_check;


// 变量节点121的接口
wire [17:0] value_check_to_variable_121;
wire [2:0] enable_check_to_variable_121;
wire [5:0] value_variable_121_to_decision;
wire [17:0] value_variable_121_to_check;

wire enable_variable_121_to_check;
// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_121[5:0] = value_check_53_to_variable_121;
assign enable_check_to_variable_121[0] = enable_check_53_to_variable_121;
// 将变量节点121的输出与校验节点53的输入相连
assign value_variable_121_to_check_53 = value_variable_121_to_check[5:0];
assign enable_variable_121_to_check_53 = enable_variable_121_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_121[11:6] = value_check_91_to_variable_121;
assign enable_check_to_variable_121[1] = enable_check_91_to_variable_121;
// 将变量节点121的输出与校验节点91的输入相连
assign value_variable_121_to_check_91 = value_variable_121_to_check[11:6];
assign enable_variable_121_to_check_91 = enable_variable_121_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_121[17:12] = value_check_116_to_variable_121;
assign enable_check_to_variable_121[2] = enable_check_116_to_variable_121;
// 将变量节点121的输出与校验节点116的输入相连
assign value_variable_121_to_check_116 = value_variable_121_to_check[17:12];
assign enable_variable_121_to_check_116 = enable_variable_121_to_check;


// 变量节点122的接口
wire [17:0] value_check_to_variable_122;
wire [2:0] enable_check_to_variable_122;
wire [5:0] value_variable_122_to_decision;
wire [17:0] value_variable_122_to_check;

wire enable_variable_122_to_check;
// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_122[5:0] = value_check_60_to_variable_122;
assign enable_check_to_variable_122[0] = enable_check_60_to_variable_122;
// 将变量节点122的输出与校验节点60的输入相连
assign value_variable_122_to_check_60 = value_variable_122_to_check[5:0];
assign enable_variable_122_to_check_60 = enable_variable_122_to_check;

// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_122[11:6] = value_check_80_to_variable_122;
assign enable_check_to_variable_122[1] = enable_check_80_to_variable_122;
// 将变量节点122的输出与校验节点80的输入相连
assign value_variable_122_to_check_80 = value_variable_122_to_check[11:6];
assign enable_variable_122_to_check_80 = enable_variable_122_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_122[17:12] = value_check_89_to_variable_122;
assign enable_check_to_variable_122[2] = enable_check_89_to_variable_122;
// 将变量节点122的输出与校验节点89的输入相连
assign value_variable_122_to_check_89 = value_variable_122_to_check[17:12];
assign enable_variable_122_to_check_89 = enable_variable_122_to_check;


// 变量节点123的接口
wire [17:0] value_check_to_variable_123;
wire [2:0] enable_check_to_variable_123;
wire [5:0] value_variable_123_to_decision;
wire [17:0] value_variable_123_to_check;

wire enable_variable_123_to_check;
// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_123[5:0] = value_check_66_to_variable_123;
assign enable_check_to_variable_123[0] = enable_check_66_to_variable_123;
// 将变量节点123的输出与校验节点66的输入相连
assign value_variable_123_to_check_66 = value_variable_123_to_check[5:0];
assign enable_variable_123_to_check_66 = enable_variable_123_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_123[11:6] = value_check_104_to_variable_123;
assign enable_check_to_variable_123[1] = enable_check_104_to_variable_123;
// 将变量节点123的输出与校验节点104的输入相连
assign value_variable_123_to_check_104 = value_variable_123_to_check[11:6];
assign enable_variable_123_to_check_104 = enable_variable_123_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_123[17:12] = value_check_115_to_variable_123;
assign enable_check_to_variable_123[2] = enable_check_115_to_variable_123;
// 将变量节点123的输出与校验节点115的输入相连
assign value_variable_123_to_check_115 = value_variable_123_to_check[17:12];
assign enable_variable_123_to_check_115 = enable_variable_123_to_check;


// 变量节点124的接口
wire [17:0] value_check_to_variable_124;
wire [2:0] enable_check_to_variable_124;
wire [5:0] value_variable_124_to_decision;
wire [17:0] value_variable_124_to_check;

wire enable_variable_124_to_check;
// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_124[5:0] = value_check_70_to_variable_124;
assign enable_check_to_variable_124[0] = enable_check_70_to_variable_124;
// 将变量节点124的输出与校验节点70的输入相连
assign value_variable_124_to_check_70 = value_variable_124_to_check[5:0];
assign enable_variable_124_to_check_70 = enable_variable_124_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_124[11:6] = value_check_81_to_variable_124;
assign enable_check_to_variable_124[1] = enable_check_81_to_variable_124;
// 将变量节点124的输出与校验节点81的输入相连
assign value_variable_124_to_check_81 = value_variable_124_to_check[11:6];
assign enable_variable_124_to_check_81 = enable_variable_124_to_check;

// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_124[17:12] = value_check_95_to_variable_124;
assign enable_check_to_variable_124[2] = enable_check_95_to_variable_124;
// 将变量节点124的输出与校验节点95的输入相连
assign value_variable_124_to_check_95 = value_variable_124_to_check[17:12];
assign enable_variable_124_to_check_95 = enable_variable_124_to_check;


// 变量节点125的接口
wire [17:0] value_check_to_variable_125;
wire [2:0] enable_check_to_variable_125;
wire [5:0] value_variable_125_to_decision;
wire [17:0] value_variable_125_to_check;

wire enable_variable_125_to_check;
// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_125[5:0] = value_check_74_to_variable_125;
assign enable_check_to_variable_125[0] = enable_check_74_to_variable_125;
// 将变量节点125的输出与校验节点74的输入相连
assign value_variable_125_to_check_74 = value_variable_125_to_check[5:0];
assign enable_variable_125_to_check_74 = enable_variable_125_to_check;

// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_125[11:6] = value_check_82_to_variable_125;
assign enable_check_to_variable_125[1] = enable_check_82_to_variable_125;
// 将变量节点125的输出与校验节点82的输入相连
assign value_variable_125_to_check_82 = value_variable_125_to_check[11:6];
assign enable_variable_125_to_check_82 = enable_variable_125_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_125[17:12] = value_check_127_to_variable_125;
assign enable_check_to_variable_125[2] = enable_check_127_to_variable_125;
// 将变量节点125的输出与校验节点127的输入相连
assign value_variable_125_to_check_127 = value_variable_125_to_check[17:12];
assign enable_variable_125_to_check_127 = enable_variable_125_to_check;


// 变量节点126的接口
wire [17:0] value_check_to_variable_126;
wire [2:0] enable_check_to_variable_126;
wire [5:0] value_variable_126_to_decision;
wire [17:0] value_variable_126_to_check;

wire enable_variable_126_to_check;
// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_126[5:0] = value_check_83_to_variable_126;
assign enable_check_to_variable_126[0] = enable_check_83_to_variable_126;
// 将变量节点126的输出与校验节点83的输入相连
assign value_variable_126_to_check_83 = value_variable_126_to_check[5:0];
assign enable_variable_126_to_check_83 = enable_variable_126_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_126[11:6] = value_check_108_to_variable_126;
assign enable_check_to_variable_126[1] = enable_check_108_to_variable_126;
// 将变量节点126的输出与校验节点108的输入相连
assign value_variable_126_to_check_108 = value_variable_126_to_check[11:6];
assign enable_variable_126_to_check_108 = enable_variable_126_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_126[17:12] = value_check_125_to_variable_126;
assign enable_check_to_variable_126[2] = enable_check_125_to_variable_126;
// 将变量节点126的输出与校验节点125的输入相连
assign value_variable_126_to_check_125 = value_variable_126_to_check[17:12];
assign enable_variable_126_to_check_125 = enable_variable_126_to_check;


// 变量节点127的接口
wire [17:0] value_check_to_variable_127;
wire [2:0] enable_check_to_variable_127;
wire [5:0] value_variable_127_to_decision;
wire [17:0] value_variable_127_to_check;

wire enable_variable_127_to_check;
// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_127[5:0] = value_check_64_to_variable_127;
assign enable_check_to_variable_127[0] = enable_check_64_to_variable_127;
// 将变量节点127的输出与校验节点64的输入相连
assign value_variable_127_to_check_64 = value_variable_127_to_check[5:0];
assign enable_variable_127_to_check_64 = enable_variable_127_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_127[11:6] = value_check_85_to_variable_127;
assign enable_check_to_variable_127[1] = enable_check_85_to_variable_127;
// 将变量节点127的输出与校验节点85的输入相连
assign value_variable_127_to_check_85 = value_variable_127_to_check[11:6];
assign enable_variable_127_to_check_85 = enable_variable_127_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_127[17:12] = value_check_106_to_variable_127;
assign enable_check_to_variable_127[2] = enable_check_106_to_variable_127;
// 将变量节点127的输出与校验节点106的输入相连
assign value_variable_127_to_check_106 = value_variable_127_to_check[17:12];
assign enable_variable_127_to_check_106 = enable_variable_127_to_check;


// 变量节点128的接口
wire [17:0] value_check_to_variable_128;
wire [2:0] enable_check_to_variable_128;
wire [5:0] value_variable_128_to_decision;
wire [17:0] value_variable_128_to_check;

wire enable_variable_128_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_128[5:0] = value_check_4_to_variable_128;
assign enable_check_to_variable_128[0] = enable_check_4_to_variable_128;
// 将变量节点128的输出与校验节点4的输入相连
assign value_variable_128_to_check_4 = value_variable_128_to_check[5:0];
assign enable_variable_128_to_check_4 = enable_variable_128_to_check;

// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_128[11:6] = value_check_86_to_variable_128;
assign enable_check_to_variable_128[1] = enable_check_86_to_variable_128;
// 将变量节点128的输出与校验节点86的输入相连
assign value_variable_128_to_check_86 = value_variable_128_to_check[11:6];
assign enable_variable_128_to_check_86 = enable_variable_128_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_128[17:12] = value_check_96_to_variable_128;
assign enable_check_to_variable_128[2] = enable_check_96_to_variable_128;
// 将变量节点128的输出与校验节点96的输入相连
assign value_variable_128_to_check_96 = value_variable_128_to_check[17:12];
assign enable_variable_128_to_check_96 = enable_variable_128_to_check;


// 变量节点129的接口
wire [17:0] value_check_to_variable_129;
wire [2:0] enable_check_to_variable_129;
wire [5:0] value_variable_129_to_decision;
wire [17:0] value_variable_129_to_check;

wire enable_variable_129_to_check;
// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_129[5:0] = value_check_37_to_variable_129;
assign enable_check_to_variable_129[0] = enable_check_37_to_variable_129;
// 将变量节点129的输出与校验节点37的输入相连
assign value_variable_129_to_check_37 = value_variable_129_to_check[5:0];
assign enable_variable_129_to_check_37 = enable_variable_129_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_129[11:6] = value_check_85_to_variable_129;
assign enable_check_to_variable_129[1] = enable_check_85_to_variable_129;
// 将变量节点129的输出与校验节点85的输入相连
assign value_variable_129_to_check_85 = value_variable_129_to_check[11:6];
assign enable_variable_129_to_check_85 = enable_variable_129_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_129[17:12] = value_check_88_to_variable_129;
assign enable_check_to_variable_129[2] = enable_check_88_to_variable_129;
// 将变量节点129的输出与校验节点88的输入相连
assign value_variable_129_to_check_88 = value_variable_129_to_check[17:12];
assign enable_variable_129_to_check_88 = enable_variable_129_to_check;


// 变量节点130的接口
wire [17:0] value_check_to_variable_130;
wire [2:0] enable_check_to_variable_130;
wire [5:0] value_variable_130_to_decision;
wire [17:0] value_variable_130_to_check;

wire enable_variable_130_to_check;
// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_130[5:0] = value_check_66_to_variable_130;
assign enable_check_to_variable_130[0] = enable_check_66_to_variable_130;
// 将变量节点130的输出与校验节点66的输入相连
assign value_variable_130_to_check_66 = value_variable_130_to_check[5:0];
assign enable_variable_130_to_check_66 = enable_variable_130_to_check;

// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_130[11:6] = value_check_74_to_variable_130;
assign enable_check_to_variable_130[1] = enable_check_74_to_variable_130;
// 将变量节点130的输出与校验节点74的输入相连
assign value_variable_130_to_check_74 = value_variable_130_to_check[11:6];
assign enable_variable_130_to_check_74 = enable_variable_130_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_130[17:12] = value_check_117_to_variable_130;
assign enable_check_to_variable_130[2] = enable_check_117_to_variable_130;
// 将变量节点130的输出与校验节点117的输入相连
assign value_variable_130_to_check_117 = value_variable_130_to_check[17:12];
assign enable_variable_130_to_check_117 = enable_variable_130_to_check;


// 变量节点131的接口
wire [17:0] value_check_to_variable_131;
wire [2:0] enable_check_to_variable_131;
wire [5:0] value_variable_131_to_decision;
wire [17:0] value_variable_131_to_check;

wire enable_variable_131_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_131[5:0] = value_check_0_to_variable_131;
assign enable_check_to_variable_131[0] = enable_check_0_to_variable_131;
// 将变量节点131的输出与校验节点0的输入相连
assign value_variable_131_to_check_0 = value_variable_131_to_check[5:0];
assign enable_variable_131_to_check_0 = enable_variable_131_to_check;

// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_131[11:6] = value_check_6_to_variable_131;
assign enable_check_to_variable_131[1] = enable_check_6_to_variable_131;
// 将变量节点131的输出与校验节点6的输入相连
assign value_variable_131_to_check_6 = value_variable_131_to_check[11:6];
assign enable_variable_131_to_check_6 = enable_variable_131_to_check;

// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_131[17:12] = value_check_76_to_variable_131;
assign enable_check_to_variable_131[2] = enable_check_76_to_variable_131;
// 将变量节点131的输出与校验节点76的输入相连
assign value_variable_131_to_check_76 = value_variable_131_to_check[17:12];
assign enable_variable_131_to_check_76 = enable_variable_131_to_check;


// 变量节点132的接口
wire [17:0] value_check_to_variable_132;
wire [2:0] enable_check_to_variable_132;
wire [5:0] value_variable_132_to_decision;
wire [17:0] value_variable_132_to_check;

wire enable_variable_132_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_132[5:0] = value_check_1_to_variable_132;
assign enable_check_to_variable_132[0] = enable_check_1_to_variable_132;
// 将变量节点132的输出与校验节点1的输入相连
assign value_variable_132_to_check_1 = value_variable_132_to_check[5:0];
assign enable_variable_132_to_check_1 = enable_variable_132_to_check;

// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_132[11:6] = value_check_21_to_variable_132;
assign enable_check_to_variable_132[1] = enable_check_21_to_variable_132;
// 将变量节点132的输出与校验节点21的输入相连
assign value_variable_132_to_check_21 = value_variable_132_to_check[11:6];
assign enable_variable_132_to_check_21 = enable_variable_132_to_check;

// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_132[17:12] = value_check_62_to_variable_132;
assign enable_check_to_variable_132[2] = enable_check_62_to_variable_132;
// 将变量节点132的输出与校验节点62的输入相连
assign value_variable_132_to_check_62 = value_variable_132_to_check[17:12];
assign enable_variable_132_to_check_62 = enable_variable_132_to_check;


// 变量节点133的接口
wire [17:0] value_check_to_variable_133;
wire [2:0] enable_check_to_variable_133;
wire [5:0] value_variable_133_to_decision;
wire [17:0] value_variable_133_to_check;

wire enable_variable_133_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_133[5:0] = value_check_2_to_variable_133;
assign enable_check_to_variable_133[0] = enable_check_2_to_variable_133;
// 将变量节点133的输出与校验节点2的输入相连
assign value_variable_133_to_check_2 = value_variable_133_to_check[5:0];
assign enable_variable_133_to_check_2 = enable_variable_133_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_133[11:6] = value_check_92_to_variable_133;
assign enable_check_to_variable_133[1] = enable_check_92_to_variable_133;
// 将变量节点133的输出与校验节点92的输入相连
assign value_variable_133_to_check_92 = value_variable_133_to_check[11:6];
assign enable_variable_133_to_check_92 = enable_variable_133_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_133[17:12] = value_check_94_to_variable_133;
assign enable_check_to_variable_133[2] = enable_check_94_to_variable_133;
// 将变量节点133的输出与校验节点94的输入相连
assign value_variable_133_to_check_94 = value_variable_133_to_check[17:12];
assign enable_variable_133_to_check_94 = enable_variable_133_to_check;


// 变量节点134的接口
wire [17:0] value_check_to_variable_134;
wire [2:0] enable_check_to_variable_134;
wire [5:0] value_variable_134_to_decision;
wire [17:0] value_variable_134_to_check;

wire enable_variable_134_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_134[5:0] = value_check_3_to_variable_134;
assign enable_check_to_variable_134[0] = enable_check_3_to_variable_134;
// 将变量节点134的输出与校验节点3的输入相连
assign value_variable_134_to_check_3 = value_variable_134_to_check[5:0];
assign enable_variable_134_to_check_3 = enable_variable_134_to_check;

// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_134[11:6] = value_check_55_to_variable_134;
assign enable_check_to_variable_134[1] = enable_check_55_to_variable_134;
// 将变量节点134的输出与校验节点55的输入相连
assign value_variable_134_to_check_55 = value_variable_134_to_check[11:6];
assign enable_variable_134_to_check_55 = enable_variable_134_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_134[17:12] = value_check_118_to_variable_134;
assign enable_check_to_variable_134[2] = enable_check_118_to_variable_134;
// 将变量节点134的输出与校验节点118的输入相连
assign value_variable_134_to_check_118 = value_variable_134_to_check[17:12];
assign enable_variable_134_to_check_118 = enable_variable_134_to_check;


// 变量节点135的接口
wire [17:0] value_check_to_variable_135;
wire [2:0] enable_check_to_variable_135;
wire [5:0] value_variable_135_to_decision;
wire [17:0] value_variable_135_to_check;

wire enable_variable_135_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_135[5:0] = value_check_5_to_variable_135;
assign enable_check_to_variable_135[0] = enable_check_5_to_variable_135;
// 将变量节点135的输出与校验节点5的输入相连
assign value_variable_135_to_check_5 = value_variable_135_to_check[5:0];
assign enable_variable_135_to_check_5 = enable_variable_135_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_135[11:6] = value_check_34_to_variable_135;
assign enable_check_to_variable_135[1] = enable_check_34_to_variable_135;
// 将变量节点135的输出与校验节点34的输入相连
assign value_variable_135_to_check_34 = value_variable_135_to_check[11:6];
assign enable_variable_135_to_check_34 = enable_variable_135_to_check;

// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_135[17:12] = value_check_35_to_variable_135;
assign enable_check_to_variable_135[2] = enable_check_35_to_variable_135;
// 将变量节点135的输出与校验节点35的输入相连
assign value_variable_135_to_check_35 = value_variable_135_to_check[17:12];
assign enable_variable_135_to_check_35 = enable_variable_135_to_check;


// 变量节点136的接口
wire [17:0] value_check_to_variable_136;
wire [2:0] enable_check_to_variable_136;
wire [5:0] value_variable_136_to_decision;
wire [17:0] value_variable_136_to_check;

wire enable_variable_136_to_check;
// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_136[5:0] = value_check_7_to_variable_136;
assign enable_check_to_variable_136[0] = enable_check_7_to_variable_136;
// 将变量节点136的输出与校验节点7的输入相连
assign value_variable_136_to_check_7 = value_variable_136_to_check[5:0];
assign enable_variable_136_to_check_7 = enable_variable_136_to_check;

// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_136[11:6] = value_check_49_to_variable_136;
assign enable_check_to_variable_136[1] = enable_check_49_to_variable_136;
// 将变量节点136的输出与校验节点49的输入相连
assign value_variable_136_to_check_49 = value_variable_136_to_check[11:6];
assign enable_variable_136_to_check_49 = enable_variable_136_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_136[17:12] = value_check_123_to_variable_136;
assign enable_check_to_variable_136[2] = enable_check_123_to_variable_136;
// 将变量节点136的输出与校验节点123的输入相连
assign value_variable_136_to_check_123 = value_variable_136_to_check[17:12];
assign enable_variable_136_to_check_123 = enable_variable_136_to_check;


// 变量节点137的接口
wire [17:0] value_check_to_variable_137;
wire [2:0] enable_check_to_variable_137;
wire [5:0] value_variable_137_to_decision;
wire [17:0] value_variable_137_to_check;

wire enable_variable_137_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_137[5:0] = value_check_8_to_variable_137;
assign enable_check_to_variable_137[0] = enable_check_8_to_variable_137;
// 将变量节点137的输出与校验节点8的输入相连
assign value_variable_137_to_check_8 = value_variable_137_to_check[5:0];
assign enable_variable_137_to_check_8 = enable_variable_137_to_check;

// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_137[11:6] = value_check_25_to_variable_137;
assign enable_check_to_variable_137[1] = enable_check_25_to_variable_137;
// 将变量节点137的输出与校验节点25的输入相连
assign value_variable_137_to_check_25 = value_variable_137_to_check[11:6];
assign enable_variable_137_to_check_25 = enable_variable_137_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_137[17:12] = value_check_90_to_variable_137;
assign enable_check_to_variable_137[2] = enable_check_90_to_variable_137;
// 将变量节点137的输出与校验节点90的输入相连
assign value_variable_137_to_check_90 = value_variable_137_to_check[17:12];
assign enable_variable_137_to_check_90 = enable_variable_137_to_check;


// 变量节点138的接口
wire [17:0] value_check_to_variable_138;
wire [2:0] enable_check_to_variable_138;
wire [5:0] value_variable_138_to_decision;
wire [17:0] value_variable_138_to_check;

wire enable_variable_138_to_check;
// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_138[5:0] = value_check_9_to_variable_138;
assign enable_check_to_variable_138[0] = enable_check_9_to_variable_138;
// 将变量节点138的输出与校验节点9的输入相连
assign value_variable_138_to_check_9 = value_variable_138_to_check[5:0];
assign enable_variable_138_to_check_9 = enable_variable_138_to_check;

// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_138[11:6] = value_check_36_to_variable_138;
assign enable_check_to_variable_138[1] = enable_check_36_to_variable_138;
// 将变量节点138的输出与校验节点36的输入相连
assign value_variable_138_to_check_36 = value_variable_138_to_check[11:6];
assign enable_variable_138_to_check_36 = enable_variable_138_to_check;

// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_138[17:12] = value_check_58_to_variable_138;
assign enable_check_to_variable_138[2] = enable_check_58_to_variable_138;
// 将变量节点138的输出与校验节点58的输入相连
assign value_variable_138_to_check_58 = value_variable_138_to_check[17:12];
assign enable_variable_138_to_check_58 = enable_variable_138_to_check;


// 变量节点139的接口
wire [17:0] value_check_to_variable_139;
wire [2:0] enable_check_to_variable_139;
wire [5:0] value_variable_139_to_decision;
wire [17:0] value_variable_139_to_check;

wire enable_variable_139_to_check;
// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_139[5:0] = value_check_10_to_variable_139;
assign enable_check_to_variable_139[0] = enable_check_10_to_variable_139;
// 将变量节点139的输出与校验节点10的输入相连
assign value_variable_139_to_check_10 = value_variable_139_to_check[5:0];
assign enable_variable_139_to_check_10 = enable_variable_139_to_check;

// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_139[11:6] = value_check_40_to_variable_139;
assign enable_check_to_variable_139[1] = enable_check_40_to_variable_139;
// 将变量节点139的输出与校验节点40的输入相连
assign value_variable_139_to_check_40 = value_variable_139_to_check[11:6];
assign enable_variable_139_to_check_40 = enable_variable_139_to_check;

// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_139[17:12] = value_check_69_to_variable_139;
assign enable_check_to_variable_139[2] = enable_check_69_to_variable_139;
// 将变量节点139的输出与校验节点69的输入相连
assign value_variable_139_to_check_69 = value_variable_139_to_check[17:12];
assign enable_variable_139_to_check_69 = enable_variable_139_to_check;


// 变量节点140的接口
wire [17:0] value_check_to_variable_140;
wire [2:0] enable_check_to_variable_140;
wire [5:0] value_variable_140_to_decision;
wire [17:0] value_variable_140_to_check;

wire enable_variable_140_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_140[5:0] = value_check_11_to_variable_140;
assign enable_check_to_variable_140[0] = enable_check_11_to_variable_140;
// 将变量节点140的输出与校验节点11的输入相连
assign value_variable_140_to_check_11 = value_variable_140_to_check[5:0];
assign enable_variable_140_to_check_11 = enable_variable_140_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_140[11:6] = value_check_77_to_variable_140;
assign enable_check_to_variable_140[1] = enable_check_77_to_variable_140;
// 将变量节点140的输出与校验节点77的输入相连
assign value_variable_140_to_check_77 = value_variable_140_to_check[11:6];
assign enable_variable_140_to_check_77 = enable_variable_140_to_check;

// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_140[17:12] = value_check_83_to_variable_140;
assign enable_check_to_variable_140[2] = enable_check_83_to_variable_140;
// 将变量节点140的输出与校验节点83的输入相连
assign value_variable_140_to_check_83 = value_variable_140_to_check[17:12];
assign enable_variable_140_to_check_83 = enable_variable_140_to_check;


// 变量节点141的接口
wire [17:0] value_check_to_variable_141;
wire [2:0] enable_check_to_variable_141;
wire [5:0] value_variable_141_to_decision;
wire [17:0] value_variable_141_to_check;

wire enable_variable_141_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_141[5:0] = value_check_13_to_variable_141;
assign enable_check_to_variable_141[0] = enable_check_13_to_variable_141;
// 将变量节点141的输出与校验节点13的输入相连
assign value_variable_141_to_check_13 = value_variable_141_to_check[5:0];
assign enable_variable_141_to_check_13 = enable_variable_141_to_check;

// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_141[11:6] = value_check_50_to_variable_141;
assign enable_check_to_variable_141[1] = enable_check_50_to_variable_141;
// 将变量节点141的输出与校验节点50的输入相连
assign value_variable_141_to_check_50 = value_variable_141_to_check[11:6];
assign enable_variable_141_to_check_50 = enable_variable_141_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_141[17:12] = value_check_75_to_variable_141;
assign enable_check_to_variable_141[2] = enable_check_75_to_variable_141;
// 将变量节点141的输出与校验节点75的输入相连
assign value_variable_141_to_check_75 = value_variable_141_to_check[17:12];
assign enable_variable_141_to_check_75 = enable_variable_141_to_check;


// 变量节点142的接口
wire [17:0] value_check_to_variable_142;
wire [2:0] enable_check_to_variable_142;
wire [5:0] value_variable_142_to_decision;
wire [17:0] value_variable_142_to_check;

wire enable_variable_142_to_check;
// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_142[5:0] = value_check_14_to_variable_142;
assign enable_check_to_variable_142[0] = enable_check_14_to_variable_142;
// 将变量节点142的输出与校验节点14的输入相连
assign value_variable_142_to_check_14 = value_variable_142_to_check[5:0];
assign enable_variable_142_to_check_14 = enable_variable_142_to_check;

// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_142[11:6] = value_check_41_to_variable_142;
assign enable_check_to_variable_142[1] = enable_check_41_to_variable_142;
// 将变量节点142的输出与校验节点41的输入相连
assign value_variable_142_to_check_41 = value_variable_142_to_check[11:6];
assign enable_variable_142_to_check_41 = enable_variable_142_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_142[17:12] = value_check_117_to_variable_142;
assign enable_check_to_variable_142[2] = enable_check_117_to_variable_142;
// 将变量节点142的输出与校验节点117的输入相连
assign value_variable_142_to_check_117 = value_variable_142_to_check[17:12];
assign enable_variable_142_to_check_117 = enable_variable_142_to_check;


// 变量节点143的接口
wire [17:0] value_check_to_variable_143;
wire [2:0] enable_check_to_variable_143;
wire [5:0] value_variable_143_to_decision;
wire [17:0] value_variable_143_to_check;

wire enable_variable_143_to_check;
// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_143[5:0] = value_check_15_to_variable_143;
assign enable_check_to_variable_143[0] = enable_check_15_to_variable_143;
// 将变量节点143的输出与校验节点15的输入相连
assign value_variable_143_to_check_15 = value_variable_143_to_check[5:0];
assign enable_variable_143_to_check_15 = enable_variable_143_to_check;

// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_143[11:6] = value_check_43_to_variable_143;
assign enable_check_to_variable_143[1] = enable_check_43_to_variable_143;
// 将变量节点143的输出与校验节点43的输入相连
assign value_variable_143_to_check_43 = value_variable_143_to_check[11:6];
assign enable_variable_143_to_check_43 = enable_variable_143_to_check;

// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_143[17:12] = value_check_47_to_variable_143;
assign enable_check_to_variable_143[2] = enable_check_47_to_variable_143;
// 将变量节点143的输出与校验节点47的输入相连
assign value_variable_143_to_check_47 = value_variable_143_to_check[17:12];
assign enable_variable_143_to_check_47 = enable_variable_143_to_check;


// 变量节点144的接口
wire [17:0] value_check_to_variable_144;
wire [2:0] enable_check_to_variable_144;
wire [5:0] value_variable_144_to_decision;
wire [17:0] value_variable_144_to_check;

wire enable_variable_144_to_check;
// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_144[5:0] = value_check_16_to_variable_144;
assign enable_check_to_variable_144[0] = enable_check_16_to_variable_144;
// 将变量节点144的输出与校验节点16的输入相连
assign value_variable_144_to_check_16 = value_variable_144_to_check[5:0];
assign enable_variable_144_to_check_16 = enable_variable_144_to_check;

// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_144[11:6] = value_check_42_to_variable_144;
assign enable_check_to_variable_144[1] = enable_check_42_to_variable_144;
// 将变量节点144的输出与校验节点42的输入相连
assign value_variable_144_to_check_42 = value_variable_144_to_check[11:6];
assign enable_variable_144_to_check_42 = enable_variable_144_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_144[17:12] = value_check_104_to_variable_144;
assign enable_check_to_variable_144[2] = enable_check_104_to_variable_144;
// 将变量节点144的输出与校验节点104的输入相连
assign value_variable_144_to_check_104 = value_variable_144_to_check[17:12];
assign enable_variable_144_to_check_104 = enable_variable_144_to_check;


// 变量节点145的接口
wire [17:0] value_check_to_variable_145;
wire [2:0] enable_check_to_variable_145;
wire [5:0] value_variable_145_to_decision;
wire [17:0] value_variable_145_to_check;

wire enable_variable_145_to_check;
// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_145[5:0] = value_check_17_to_variable_145;
assign enable_check_to_variable_145[0] = enable_check_17_to_variable_145;
// 将变量节点145的输出与校验节点17的输入相连
assign value_variable_145_to_check_17 = value_variable_145_to_check[5:0];
assign enable_variable_145_to_check_17 = enable_variable_145_to_check;

// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_145[11:6] = value_check_18_to_variable_145;
assign enable_check_to_variable_145[1] = enable_check_18_to_variable_145;
// 将变量节点145的输出与校验节点18的输入相连
assign value_variable_145_to_check_18 = value_variable_145_to_check[11:6];
assign enable_variable_145_to_check_18 = enable_variable_145_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_145[17:12] = value_check_112_to_variable_145;
assign enable_check_to_variable_145[2] = enable_check_112_to_variable_145;
// 将变量节点145的输出与校验节点112的输入相连
assign value_variable_145_to_check_112 = value_variable_145_to_check[17:12];
assign enable_variable_145_to_check_112 = enable_variable_145_to_check;


// 变量节点146的接口
wire [17:0] value_check_to_variable_146;
wire [2:0] enable_check_to_variable_146;
wire [5:0] value_variable_146_to_decision;
wire [17:0] value_variable_146_to_check;

wire enable_variable_146_to_check;
// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_146[5:0] = value_check_19_to_variable_146;
assign enable_check_to_variable_146[0] = enable_check_19_to_variable_146;
// 将变量节点146的输出与校验节点19的输入相连
assign value_variable_146_to_check_19 = value_variable_146_to_check[5:0];
assign enable_variable_146_to_check_19 = enable_variable_146_to_check;

// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_146[11:6] = value_check_39_to_variable_146;
assign enable_check_to_variable_146[1] = enable_check_39_to_variable_146;
// 将变量节点146的输出与校验节点39的输入相连
assign value_variable_146_to_check_39 = value_variable_146_to_check[11:6];
assign enable_variable_146_to_check_39 = enable_variable_146_to_check;

// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_146[17:12] = value_check_59_to_variable_146;
assign enable_check_to_variable_146[2] = enable_check_59_to_variable_146;
// 将变量节点146的输出与校验节点59的输入相连
assign value_variable_146_to_check_59 = value_variable_146_to_check[17:12];
assign enable_variable_146_to_check_59 = enable_variable_146_to_check;


// 变量节点147的接口
wire [17:0] value_check_to_variable_147;
wire [2:0] enable_check_to_variable_147;
wire [5:0] value_variable_147_to_decision;
wire [17:0] value_variable_147_to_check;

wire enable_variable_147_to_check;
// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_147[5:0] = value_check_20_to_variable_147;
assign enable_check_to_variable_147[0] = enable_check_20_to_variable_147;
// 将变量节点147的输出与校验节点20的输入相连
assign value_variable_147_to_check_20 = value_variable_147_to_check[5:0];
assign enable_variable_147_to_check_20 = enable_variable_147_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_147[11:6] = value_check_89_to_variable_147;
assign enable_check_to_variable_147[1] = enable_check_89_to_variable_147;
// 将变量节点147的输出与校验节点89的输入相连
assign value_variable_147_to_check_89 = value_variable_147_to_check[11:6];
assign enable_variable_147_to_check_89 = enable_variable_147_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_147[17:12] = value_check_122_to_variable_147;
assign enable_check_to_variable_147[2] = enable_check_122_to_variable_147;
// 将变量节点147的输出与校验节点122的输入相连
assign value_variable_147_to_check_122 = value_variable_147_to_check[17:12];
assign enable_variable_147_to_check_122 = enable_variable_147_to_check;


// 变量节点148的接口
wire [17:0] value_check_to_variable_148;
wire [2:0] enable_check_to_variable_148;
wire [5:0] value_variable_148_to_decision;
wire [17:0] value_variable_148_to_check;

wire enable_variable_148_to_check;
// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_148[5:0] = value_check_22_to_variable_148;
assign enable_check_to_variable_148[0] = enable_check_22_to_variable_148;
// 将变量节点148的输出与校验节点22的输入相连
assign value_variable_148_to_check_22 = value_variable_148_to_check[5:0];
assign enable_variable_148_to_check_22 = enable_variable_148_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_148[11:6] = value_check_81_to_variable_148;
assign enable_check_to_variable_148[1] = enable_check_81_to_variable_148;
// 将变量节点148的输出与校验节点81的输入相连
assign value_variable_148_to_check_81 = value_variable_148_to_check[11:6];
assign enable_variable_148_to_check_81 = enable_variable_148_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_148[17:12] = value_check_102_to_variable_148;
assign enable_check_to_variable_148[2] = enable_check_102_to_variable_148;
// 将变量节点148的输出与校验节点102的输入相连
assign value_variable_148_to_check_102 = value_variable_148_to_check[17:12];
assign enable_variable_148_to_check_102 = enable_variable_148_to_check;


// 变量节点149的接口
wire [17:0] value_check_to_variable_149;
wire [2:0] enable_check_to_variable_149;
wire [5:0] value_variable_149_to_decision;
wire [17:0] value_variable_149_to_check;

wire enable_variable_149_to_check;
// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_149[5:0] = value_check_23_to_variable_149;
assign enable_check_to_variable_149[0] = enable_check_23_to_variable_149;
// 将变量节点149的输出与校验节点23的输入相连
assign value_variable_149_to_check_23 = value_variable_149_to_check[5:0];
assign enable_variable_149_to_check_23 = enable_variable_149_to_check;

// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_149[11:6] = value_check_60_to_variable_149;
assign enable_check_to_variable_149[1] = enable_check_60_to_variable_149;
// 将变量节点149的输出与校验节点60的输入相连
assign value_variable_149_to_check_60 = value_variable_149_to_check[11:6];
assign enable_variable_149_to_check_60 = enable_variable_149_to_check;

// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_149[17:12] = value_check_97_to_variable_149;
assign enable_check_to_variable_149[2] = enable_check_97_to_variable_149;
// 将变量节点149的输出与校验节点97的输入相连
assign value_variable_149_to_check_97 = value_variable_149_to_check[17:12];
assign enable_variable_149_to_check_97 = enable_variable_149_to_check;


// 变量节点150的接口
wire [17:0] value_check_to_variable_150;
wire [2:0] enable_check_to_variable_150;
wire [5:0] value_variable_150_to_decision;
wire [17:0] value_variable_150_to_check;

wire enable_variable_150_to_check;
// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_150[5:0] = value_check_24_to_variable_150;
assign enable_check_to_variable_150[0] = enable_check_24_to_variable_150;
// 将变量节点150的输出与校验节点24的输入相连
assign value_variable_150_to_check_24 = value_variable_150_to_check[5:0];
assign enable_variable_150_to_check_24 = enable_variable_150_to_check;

// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_150[11:6] = value_check_51_to_variable_150;
assign enable_check_to_variable_150[1] = enable_check_51_to_variable_150;
// 将变量节点150的输出与校验节点51的输入相连
assign value_variable_150_to_check_51 = value_variable_150_to_check[11:6];
assign enable_variable_150_to_check_51 = enable_variable_150_to_check;

// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_150[17:12] = value_check_70_to_variable_150;
assign enable_check_to_variable_150[2] = enable_check_70_to_variable_150;
// 将变量节点150的输出与校验节点70的输入相连
assign value_variable_150_to_check_70 = value_variable_150_to_check[17:12];
assign enable_variable_150_to_check_70 = enable_variable_150_to_check;


// 变量节点151的接口
wire [17:0] value_check_to_variable_151;
wire [2:0] enable_check_to_variable_151;
wire [5:0] value_variable_151_to_decision;
wire [17:0] value_variable_151_to_check;

wire enable_variable_151_to_check;
// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_151[5:0] = value_check_26_to_variable_151;
assign enable_check_to_variable_151[0] = enable_check_26_to_variable_151;
// 将变量节点151的输出与校验节点26的输入相连
assign value_variable_151_to_check_26 = value_variable_151_to_check[5:0];
assign enable_variable_151_to_check_26 = enable_variable_151_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_151[11:6] = value_check_61_to_variable_151;
assign enable_check_to_variable_151[1] = enable_check_61_to_variable_151;
// 将变量节点151的输出与校验节点61的输入相连
assign value_variable_151_to_check_61 = value_variable_151_to_check[11:6];
assign enable_variable_151_to_check_61 = enable_variable_151_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_151[17:12] = value_check_96_to_variable_151;
assign enable_check_to_variable_151[2] = enable_check_96_to_variable_151;
// 将变量节点151的输出与校验节点96的输入相连
assign value_variable_151_to_check_96 = value_variable_151_to_check[17:12];
assign enable_variable_151_to_check_96 = enable_variable_151_to_check;


// 变量节点152的接口
wire [17:0] value_check_to_variable_152;
wire [2:0] enable_check_to_variable_152;
wire [5:0] value_variable_152_to_decision;
wire [17:0] value_variable_152_to_check;

wire enable_variable_152_to_check;
// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_152[5:0] = value_check_27_to_variable_152;
assign enable_check_to_variable_152[0] = enable_check_27_to_variable_152;
// 将变量节点152的输出与校验节点27的输入相连
assign value_variable_152_to_check_27 = value_variable_152_to_check[5:0];
assign enable_variable_152_to_check_27 = enable_variable_152_to_check;

// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_152[11:6] = value_check_53_to_variable_152;
assign enable_check_to_variable_152[1] = enable_check_53_to_variable_152;
// 将变量节点152的输出与校验节点53的输入相连
assign value_variable_152_to_check_53 = value_variable_152_to_check[11:6];
assign enable_variable_152_to_check_53 = enable_variable_152_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_152[17:12] = value_check_118_to_variable_152;
assign enable_check_to_variable_152[2] = enable_check_118_to_variable_152;
// 将变量节点152的输出与校验节点118的输入相连
assign value_variable_152_to_check_118 = value_variable_152_to_check[17:12];
assign enable_variable_152_to_check_118 = enable_variable_152_to_check;


// 变量节点153的接口
wire [17:0] value_check_to_variable_153;
wire [2:0] enable_check_to_variable_153;
wire [5:0] value_variable_153_to_decision;
wire [17:0] value_variable_153_to_check;

wire enable_variable_153_to_check;
// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_153[5:0] = value_check_28_to_variable_153;
assign enable_check_to_variable_153[0] = enable_check_28_to_variable_153;
// 将变量节点153的输出与校验节点28的输入相连
assign value_variable_153_to_check_28 = value_variable_153_to_check[5:0];
assign enable_variable_153_to_check_28 = enable_variable_153_to_check;

// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_153[11:6] = value_check_46_to_variable_153;
assign enable_check_to_variable_153[1] = enable_check_46_to_variable_153;
// 将变量节点153的输出与校验节点46的输入相连
assign value_variable_153_to_check_46 = value_variable_153_to_check[11:6];
assign enable_variable_153_to_check_46 = enable_variable_153_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_153[17:12] = value_check_111_to_variable_153;
assign enable_check_to_variable_153[2] = enable_check_111_to_variable_153;
// 将变量节点153的输出与校验节点111的输入相连
assign value_variable_153_to_check_111 = value_variable_153_to_check[17:12];
assign enable_variable_153_to_check_111 = enable_variable_153_to_check;


// 变量节点154的接口
wire [17:0] value_check_to_variable_154;
wire [2:0] enable_check_to_variable_154;
wire [5:0] value_variable_154_to_decision;
wire [17:0] value_variable_154_to_check;

wire enable_variable_154_to_check;
// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_154[5:0] = value_check_29_to_variable_154;
assign enable_check_to_variable_154[0] = enable_check_29_to_variable_154;
// 将变量节点154的输出与校验节点29的输入相连
assign value_variable_154_to_check_29 = value_variable_154_to_check[5:0];
assign enable_variable_154_to_check_29 = enable_variable_154_to_check;

// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_154[11:6] = value_check_109_to_variable_154;
assign enable_check_to_variable_154[1] = enable_check_109_to_variable_154;
// 将变量节点154的输出与校验节点109的输入相连
assign value_variable_154_to_check_109 = value_variable_154_to_check[11:6];
assign enable_variable_154_to_check_109 = enable_variable_154_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_154[17:12] = value_check_126_to_variable_154;
assign enable_check_to_variable_154[2] = enable_check_126_to_variable_154;
// 将变量节点154的输出与校验节点126的输入相连
assign value_variable_154_to_check_126 = value_variable_154_to_check[17:12];
assign enable_variable_154_to_check_126 = enable_variable_154_to_check;


// 变量节点155的接口
wire [17:0] value_check_to_variable_155;
wire [2:0] enable_check_to_variable_155;
wire [5:0] value_variable_155_to_decision;
wire [17:0] value_variable_155_to_check;

wire enable_variable_155_to_check;
// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_155[5:0] = value_check_30_to_variable_155;
assign enable_check_to_variable_155[0] = enable_check_30_to_variable_155;
// 将变量节点155的输出与校验节点30的输入相连
assign value_variable_155_to_check_30 = value_variable_155_to_check[5:0];
assign enable_variable_155_to_check_30 = enable_variable_155_to_check;

// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_155[11:6] = value_check_38_to_variable_155;
assign enable_check_to_variable_155[1] = enable_check_38_to_variable_155;
// 将变量节点155的输出与校验节点38的输入相连
assign value_variable_155_to_check_38 = value_variable_155_to_check[11:6];
assign enable_variable_155_to_check_38 = enable_variable_155_to_check;

// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_155[17:12] = value_check_80_to_variable_155;
assign enable_check_to_variable_155[2] = enable_check_80_to_variable_155;
// 将变量节点155的输出与校验节点80的输入相连
assign value_variable_155_to_check_80 = value_variable_155_to_check[17:12];
assign enable_variable_155_to_check_80 = enable_variable_155_to_check;


// 变量节点156的接口
wire [17:0] value_check_to_variable_156;
wire [2:0] enable_check_to_variable_156;
wire [5:0] value_variable_156_to_decision;
wire [17:0] value_variable_156_to_check;

wire enable_variable_156_to_check;
// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_156[5:0] = value_check_31_to_variable_156;
assign enable_check_to_variable_156[0] = enable_check_31_to_variable_156;
// 将变量节点156的输出与校验节点31的输入相连
assign value_variable_156_to_check_31 = value_variable_156_to_check[5:0];
assign enable_variable_156_to_check_31 = enable_variable_156_to_check;

// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_156[11:6] = value_check_63_to_variable_156;
assign enable_check_to_variable_156[1] = enable_check_63_to_variable_156;
// 将变量节点156的输出与校验节点63的输入相连
assign value_variable_156_to_check_63 = value_variable_156_to_check[11:6];
assign enable_variable_156_to_check_63 = enable_variable_156_to_check;

// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_156[17:12] = value_check_73_to_variable_156;
assign enable_check_to_variable_156[2] = enable_check_73_to_variable_156;
// 将变量节点156的输出与校验节点73的输入相连
assign value_variable_156_to_check_73 = value_variable_156_to_check[17:12];
assign enable_variable_156_to_check_73 = enable_variable_156_to_check;


// 变量节点157的接口
wire [17:0] value_check_to_variable_157;
wire [2:0] enable_check_to_variable_157;
wire [5:0] value_variable_157_to_decision;
wire [17:0] value_variable_157_to_check;

wire enable_variable_157_to_check;
// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_157[5:0] = value_check_32_to_variable_157;
assign enable_check_to_variable_157[0] = enable_check_32_to_variable_157;
// 将变量节点157的输出与校验节点32的输入相连
assign value_variable_157_to_check_32 = value_variable_157_to_check[5:0];
assign enable_variable_157_to_check_32 = enable_variable_157_to_check;

// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_157[11:6] = value_check_44_to_variable_157;
assign enable_check_to_variable_157[1] = enable_check_44_to_variable_157;
// 将变量节点157的输出与校验节点44的输入相连
assign value_variable_157_to_check_44 = value_variable_157_to_check[11:6];
assign enable_variable_157_to_check_44 = enable_variable_157_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_157[17:12] = value_check_120_to_variable_157;
assign enable_check_to_variable_157[2] = enable_check_120_to_variable_157;
// 将变量节点157的输出与校验节点120的输入相连
assign value_variable_157_to_check_120 = value_variable_157_to_check[17:12];
assign enable_variable_157_to_check_120 = enable_variable_157_to_check;


// 变量节点158的接口
wire [17:0] value_check_to_variable_158;
wire [2:0] enable_check_to_variable_158;
wire [5:0] value_variable_158_to_decision;
wire [17:0] value_variable_158_to_check;

wire enable_variable_158_to_check;
// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_158[5:0] = value_check_33_to_variable_158;
assign enable_check_to_variable_158[0] = enable_check_33_to_variable_158;
// 将变量节点158的输出与校验节点33的输入相连
assign value_variable_158_to_check_33 = value_variable_158_to_check[5:0];
assign enable_variable_158_to_check_33 = enable_variable_158_to_check;

// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_158[11:6] = value_check_71_to_variable_158;
assign enable_check_to_variable_158[1] = enable_check_71_to_variable_158;
// 将变量节点158的输出与校验节点71的输入相连
assign value_variable_158_to_check_71 = value_variable_158_to_check[11:6];
assign enable_variable_158_to_check_71 = enable_variable_158_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_158[17:12] = value_check_101_to_variable_158;
assign enable_check_to_variable_158[2] = enable_check_101_to_variable_158;
// 将变量节点158的输出与校验节点101的输入相连
assign value_variable_158_to_check_101 = value_variable_158_to_check[17:12];
assign enable_variable_158_to_check_101 = enable_variable_158_to_check;


// 变量节点159的接口
wire [17:0] value_check_to_variable_159;
wire [2:0] enable_check_to_variable_159;
wire [5:0] value_variable_159_to_decision;
wire [17:0] value_variable_159_to_check;

wire enable_variable_159_to_check;
// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_159[5:0] = value_check_45_to_variable_159;
assign enable_check_to_variable_159[0] = enable_check_45_to_variable_159;
// 将变量节点159的输出与校验节点45的输入相连
assign value_variable_159_to_check_45 = value_variable_159_to_check[5:0];
assign enable_variable_159_to_check_45 = enable_variable_159_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_159[11:6] = value_check_84_to_variable_159;
assign enable_check_to_variable_159[1] = enable_check_84_to_variable_159;
// 将变量节点159的输出与校验节点84的输入相连
assign value_variable_159_to_check_84 = value_variable_159_to_check[11:6];
assign enable_variable_159_to_check_84 = enable_variable_159_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_159[17:12] = value_check_115_to_variable_159;
assign enable_check_to_variable_159[2] = enable_check_115_to_variable_159;
// 将变量节点159的输出与校验节点115的输入相连
assign value_variable_159_to_check_115 = value_variable_159_to_check[17:12];
assign enable_variable_159_to_check_115 = enable_variable_159_to_check;


// 变量节点160的接口
wire [17:0] value_check_to_variable_160;
wire [2:0] enable_check_to_variable_160;
wire [5:0] value_variable_160_to_decision;
wire [17:0] value_variable_160_to_check;

wire enable_variable_160_to_check;
// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_160[5:0] = value_check_48_to_variable_160;
assign enable_check_to_variable_160[0] = enable_check_48_to_variable_160;
// 将变量节点160的输出与校验节点48的输入相连
assign value_variable_160_to_check_48 = value_variable_160_to_check[5:0];
assign enable_variable_160_to_check_48 = enable_variable_160_to_check;

// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_160[11:6] = value_check_65_to_variable_160;
assign enable_check_to_variable_160[1] = enable_check_65_to_variable_160;
// 将变量节点160的输出与校验节点65的输入相连
assign value_variable_160_to_check_65 = value_variable_160_to_check[11:6];
assign enable_variable_160_to_check_65 = enable_variable_160_to_check;

// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_160[17:12] = value_check_68_to_variable_160;
assign enable_check_to_variable_160[2] = enable_check_68_to_variable_160;
// 将变量节点160的输出与校验节点68的输入相连
assign value_variable_160_to_check_68 = value_variable_160_to_check[17:12];
assign enable_variable_160_to_check_68 = enable_variable_160_to_check;


// 变量节点161的接口
wire [17:0] value_check_to_variable_161;
wire [2:0] enable_check_to_variable_161;
wire [5:0] value_variable_161_to_decision;
wire [17:0] value_variable_161_to_check;

wire enable_variable_161_to_check;
// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_161[5:0] = value_check_52_to_variable_161;
assign enable_check_to_variable_161[0] = enable_check_52_to_variable_161;
// 将变量节点161的输出与校验节点52的输入相连
assign value_variable_161_to_check_52 = value_variable_161_to_check[5:0];
assign enable_variable_161_to_check_52 = enable_variable_161_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_161[11:6] = value_check_91_to_variable_161;
assign enable_check_to_variable_161[1] = enable_check_91_to_variable_161;
// 将变量节点161的输出与校验节点91的输入相连
assign value_variable_161_to_check_91 = value_variable_161_to_check[11:6];
assign enable_variable_161_to_check_91 = enable_variable_161_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_161[17:12] = value_check_93_to_variable_161;
assign enable_check_to_variable_161[2] = enable_check_93_to_variable_161;
// 将变量节点161的输出与校验节点93的输入相连
assign value_variable_161_to_check_93 = value_variable_161_to_check[17:12];
assign enable_variable_161_to_check_93 = enable_variable_161_to_check;


// 变量节点162的接口
wire [17:0] value_check_to_variable_162;
wire [2:0] enable_check_to_variable_162;
wire [5:0] value_variable_162_to_decision;
wire [17:0] value_variable_162_to_check;

wire enable_variable_162_to_check;
// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_162[5:0] = value_check_54_to_variable_162;
assign enable_check_to_variable_162[0] = enable_check_54_to_variable_162;
// 将变量节点162的输出与校验节点54的输入相连
assign value_variable_162_to_check_54 = value_variable_162_to_check[5:0];
assign enable_variable_162_to_check_54 = enable_variable_162_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_162[11:6] = value_check_87_to_variable_162;
assign enable_check_to_variable_162[1] = enable_check_87_to_variable_162;
// 将变量节点162的输出与校验节点87的输入相连
assign value_variable_162_to_check_87 = value_variable_162_to_check[11:6];
assign enable_variable_162_to_check_87 = enable_variable_162_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_162[17:12] = value_check_107_to_variable_162;
assign enable_check_to_variable_162[2] = enable_check_107_to_variable_162;
// 将变量节点162的输出与校验节点107的输入相连
assign value_variable_162_to_check_107 = value_variable_162_to_check[17:12];
assign enable_variable_162_to_check_107 = enable_variable_162_to_check;


// 变量节点163的接口
wire [17:0] value_check_to_variable_163;
wire [2:0] enable_check_to_variable_163;
wire [5:0] value_variable_163_to_decision;
wire [17:0] value_variable_163_to_check;

wire enable_variable_163_to_check;
// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_163[5:0] = value_check_56_to_variable_163;
assign enable_check_to_variable_163[0] = enable_check_56_to_variable_163;
// 将变量节点163的输出与校验节点56的输入相连
assign value_variable_163_to_check_56 = value_variable_163_to_check[5:0];
assign enable_variable_163_to_check_56 = enable_variable_163_to_check;

// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_163[11:6] = value_check_79_to_variable_163;
assign enable_check_to_variable_163[1] = enable_check_79_to_variable_163;
// 将变量节点163的输出与校验节点79的输入相连
assign value_variable_163_to_check_79 = value_variable_163_to_check[11:6];
assign enable_variable_163_to_check_79 = enable_variable_163_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_163[17:12] = value_check_113_to_variable_163;
assign enable_check_to_variable_163[2] = enable_check_113_to_variable_163;
// 将变量节点163的输出与校验节点113的输入相连
assign value_variable_163_to_check_113 = value_variable_163_to_check[17:12];
assign enable_variable_163_to_check_113 = enable_variable_163_to_check;


// 变量节点164的接口
wire [17:0] value_check_to_variable_164;
wire [2:0] enable_check_to_variable_164;
wire [5:0] value_variable_164_to_decision;
wire [17:0] value_variable_164_to_check;

wire enable_variable_164_to_check;
// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_164[5:0] = value_check_64_to_variable_164;
assign enable_check_to_variable_164[0] = enable_check_64_to_variable_164;
// 将变量节点164的输出与校验节点64的输入相连
assign value_variable_164_to_check_64 = value_variable_164_to_check[5:0];
assign enable_variable_164_to_check_64 = enable_variable_164_to_check;

// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_164[11:6] = value_check_67_to_variable_164;
assign enable_check_to_variable_164[1] = enable_check_67_to_variable_164;
// 将变量节点164的输出与校验节点67的输入相连
assign value_variable_164_to_check_67 = value_variable_164_to_check[11:6];
assign enable_variable_164_to_check_67 = enable_variable_164_to_check;

// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_164[17:12] = value_check_82_to_variable_164;
assign enable_check_to_variable_164[2] = enable_check_82_to_variable_164;
// 将变量节点164的输出与校验节点82的输入相连
assign value_variable_164_to_check_82 = value_variable_164_to_check[17:12];
assign enable_variable_164_to_check_82 = enable_variable_164_to_check;


// 变量节点165的接口
wire [17:0] value_check_to_variable_165;
wire [2:0] enable_check_to_variable_165;
wire [5:0] value_variable_165_to_decision;
wire [17:0] value_variable_165_to_check;

wire enable_variable_165_to_check;
// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_165[5:0] = value_check_20_to_variable_165;
assign enable_check_to_variable_165[0] = enable_check_20_to_variable_165;
// 将变量节点165的输出与校验节点20的输入相连
assign value_variable_165_to_check_20 = value_variable_165_to_check[5:0];
assign enable_variable_165_to_check_20 = enable_variable_165_to_check;

// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_165[11:6] = value_check_72_to_variable_165;
assign enable_check_to_variable_165[1] = enable_check_72_to_variable_165;
// 将变量节点165的输出与校验节点72的输入相连
assign value_variable_165_to_check_72 = value_variable_165_to_check[11:6];
assign enable_variable_165_to_check_72 = enable_variable_165_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_165[17:12] = value_check_103_to_variable_165;
assign enable_check_to_variable_165[2] = enable_check_103_to_variable_165;
// 将变量节点165的输出与校验节点103的输入相连
assign value_variable_165_to_check_103 = value_variable_165_to_check[17:12];
assign enable_variable_165_to_check_103 = enable_variable_165_to_check;


// 变量节点166的接口
wire [17:0] value_check_to_variable_166;
wire [2:0] enable_check_to_variable_166;
wire [5:0] value_variable_166_to_decision;
wire [17:0] value_variable_166_to_check;

wire enable_variable_166_to_check;
// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_166[5:0] = value_check_86_to_variable_166;
assign enable_check_to_variable_166[0] = enable_check_86_to_variable_166;
// 将变量节点166的输出与校验节点86的输入相连
assign value_variable_166_to_check_86 = value_variable_166_to_check[5:0];
assign enable_variable_166_to_check_86 = enable_variable_166_to_check;

// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_166[11:6] = value_check_100_to_variable_166;
assign enable_check_to_variable_166[1] = enable_check_100_to_variable_166;
// 将变量节点166的输出与校验节点100的输入相连
assign value_variable_166_to_check_100 = value_variable_166_to_check[11:6];
assign enable_variable_166_to_check_100 = enable_variable_166_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_166[17:12] = value_check_106_to_variable_166;
assign enable_check_to_variable_166[2] = enable_check_106_to_variable_166;
// 将变量节点166的输出与校验节点106的输入相连
assign value_variable_166_to_check_106 = value_variable_166_to_check[17:12];
assign enable_variable_166_to_check_106 = enable_variable_166_to_check;


// 变量节点167的接口
wire [17:0] value_check_to_variable_167;
wire [2:0] enable_check_to_variable_167;
wire [5:0] value_variable_167_to_decision;
wire [17:0] value_variable_167_to_check;

wire enable_variable_167_to_check;
// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_167[5:0] = value_check_50_to_variable_167;
assign enable_check_to_variable_167[0] = enable_check_50_to_variable_167;
// 将变量节点167的输出与校验节点50的输入相连
assign value_variable_167_to_check_50 = value_variable_167_to_check[5:0];
assign enable_variable_167_to_check_50 = enable_variable_167_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_167[11:6] = value_check_88_to_variable_167;
assign enable_check_to_variable_167[1] = enable_check_88_to_variable_167;
// 将变量节点167的输出与校验节点88的输入相连
assign value_variable_167_to_check_88 = value_variable_167_to_check[11:6];
assign enable_variable_167_to_check_88 = enable_variable_167_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_167[17:12] = value_check_124_to_variable_167;
assign enable_check_to_variable_167[2] = enable_check_124_to_variable_167;
// 将变量节点167的输出与校验节点124的输入相连
assign value_variable_167_to_check_124 = value_variable_167_to_check[17:12];
assign enable_variable_167_to_check_124 = enable_variable_167_to_check;


// 变量节点168的接口
wire [17:0] value_check_to_variable_168;
wire [2:0] enable_check_to_variable_168;
wire [5:0] value_variable_168_to_decision;
wire [17:0] value_variable_168_to_check;

wire enable_variable_168_to_check;
// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_168[5:0] = value_check_95_to_variable_168;
assign enable_check_to_variable_168[0] = enable_check_95_to_variable_168;
// 将变量节点168的输出与校验节点95的输入相连
assign value_variable_168_to_check_95 = value_variable_168_to_check[5:0];
assign enable_variable_168_to_check_95 = enable_variable_168_to_check;

// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_168[11:6] = value_check_99_to_variable_168;
assign enable_check_to_variable_168[1] = enable_check_99_to_variable_168;
// 将变量节点168的输出与校验节点99的输入相连
assign value_variable_168_to_check_99 = value_variable_168_to_check[11:6];
assign enable_variable_168_to_check_99 = enable_variable_168_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_168[17:12] = value_check_114_to_variable_168;
assign enable_check_to_variable_168[2] = enable_check_114_to_variable_168;
// 将变量节点168的输出与校验节点114的输入相连
assign value_variable_168_to_check_114 = value_variable_168_to_check[17:12];
assign enable_variable_168_to_check_114 = enable_variable_168_to_check;


// 变量节点169的接口
wire [17:0] value_check_to_variable_169;
wire [2:0] enable_check_to_variable_169;
wire [5:0] value_variable_169_to_decision;
wire [17:0] value_variable_169_to_check;

wire enable_variable_169_to_check;
// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_169[5:0] = value_check_98_to_variable_169;
assign enable_check_to_variable_169[0] = enable_check_98_to_variable_169;
// 将变量节点169的输出与校验节点98的输入相连
assign value_variable_169_to_check_98 = value_variable_169_to_check[5:0];
assign enable_variable_169_to_check_98 = enable_variable_169_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_169[11:6] = value_check_108_to_variable_169;
assign enable_check_to_variable_169[1] = enable_check_108_to_variable_169;
// 将变量节点169的输出与校验节点108的输入相连
assign value_variable_169_to_check_108 = value_variable_169_to_check[11:6];
assign enable_variable_169_to_check_108 = enable_variable_169_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_169[17:12] = value_check_121_to_variable_169;
assign enable_check_to_variable_169[2] = enable_check_121_to_variable_169;
// 将变量节点169的输出与校验节点121的输入相连
assign value_variable_169_to_check_121 = value_variable_169_to_check[17:12];
assign enable_variable_169_to_check_121 = enable_variable_169_to_check;


// 变量节点170的接口
wire [17:0] value_check_to_variable_170;
wire [2:0] enable_check_to_variable_170;
wire [5:0] value_variable_170_to_decision;
wire [17:0] value_variable_170_to_check;

wire enable_variable_170_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_170[5:0] = value_check_0_to_variable_170;
assign enable_check_to_variable_170[0] = enable_check_0_to_variable_170;
// 将变量节点170的输出与校验节点0的输入相连
assign value_variable_170_to_check_0 = value_variable_170_to_check[5:0];
assign enable_variable_170_to_check_0 = enable_variable_170_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_170[11:6] = value_check_105_to_variable_170;
assign enable_check_to_variable_170[1] = enable_check_105_to_variable_170;
// 将变量节点170的输出与校验节点105的输入相连
assign value_variable_170_to_check_105 = value_variable_170_to_check[11:6];
assign enable_variable_170_to_check_105 = enable_variable_170_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_170[17:12] = value_check_116_to_variable_170;
assign enable_check_to_variable_170[2] = enable_check_116_to_variable_170;
// 将变量节点170的输出与校验节点116的输入相连
assign value_variable_170_to_check_116 = value_variable_170_to_check[17:12];
assign enable_variable_170_to_check_116 = enable_variable_170_to_check;


// 变量节点171的接口
wire [17:0] value_check_to_variable_171;
wire [2:0] enable_check_to_variable_171;
wire [5:0] value_variable_171_to_decision;
wire [17:0] value_variable_171_to_check;

wire enable_variable_171_to_check;
// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_171[5:0] = value_check_110_to_variable_171;
assign enable_check_to_variable_171[0] = enable_check_110_to_variable_171;
// 将变量节点171的输出与校验节点110的输入相连
assign value_variable_171_to_check_110 = value_variable_171_to_check[5:0];
assign enable_variable_171_to_check_110 = enable_variable_171_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_171[11:6] = value_check_125_to_variable_171;
assign enable_check_to_variable_171[1] = enable_check_125_to_variable_171;
// 将变量节点171的输出与校验节点125的输入相连
assign value_variable_171_to_check_125 = value_variable_171_to_check[11:6];
assign enable_variable_171_to_check_125 = enable_variable_171_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_171[17:12] = value_check_127_to_variable_171;
assign enable_check_to_variable_171[2] = enable_check_127_to_variable_171;
// 将变量节点171的输出与校验节点127的输入相连
assign value_variable_171_to_check_127 = value_variable_171_to_check[17:12];
assign enable_variable_171_to_check_127 = enable_variable_171_to_check;


// 变量节点172的接口
wire [17:0] value_check_to_variable_172;
wire [2:0] enable_check_to_variable_172;
wire [5:0] value_variable_172_to_decision;
wire [17:0] value_variable_172_to_check;

wire enable_variable_172_to_check;
// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_172[5:0] = value_check_38_to_variable_172;
assign enable_check_to_variable_172[0] = enable_check_38_to_variable_172;
// 将变量节点172的输出与校验节点38的输入相连
assign value_variable_172_to_check_38 = value_variable_172_to_check[5:0];
assign enable_variable_172_to_check_38 = enable_variable_172_to_check;

// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_172[11:6] = value_check_57_to_variable_172;
assign enable_check_to_variable_172[1] = enable_check_57_to_variable_172;
// 将变量节点172的输出与校验节点57的输入相连
assign value_variable_172_to_check_57 = value_variable_172_to_check[11:6];
assign enable_variable_172_to_check_57 = enable_variable_172_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_172[17:12] = value_check_119_to_variable_172;
assign enable_check_to_variable_172[2] = enable_check_119_to_variable_172;
// 将变量节点172的输出与校验节点119的输入相连
assign value_variable_172_to_check_119 = value_variable_172_to_check[17:12];
assign enable_variable_172_to_check_119 = enable_variable_172_to_check;


// 变量节点173的接口
wire [17:0] value_check_to_variable_173;
wire [2:0] enable_check_to_variable_173;
wire [5:0] value_variable_173_to_decision;
wire [17:0] value_variable_173_to_check;

wire enable_variable_173_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_173[5:0] = value_check_1_to_variable_173;
assign enable_check_to_variable_173[0] = enable_check_1_to_variable_173;
// 将变量节点173的输出与校验节点1的输入相连
assign value_variable_173_to_check_1 = value_variable_173_to_check[5:0];
assign enable_variable_173_to_check_1 = enable_variable_173_to_check;

// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_173[11:6] = value_check_60_to_variable_173;
assign enable_check_to_variable_173[1] = enable_check_60_to_variable_173;
// 将变量节点173的输出与校验节点60的输入相连
assign value_variable_173_to_check_60 = value_variable_173_to_check[11:6];
assign enable_variable_173_to_check_60 = enable_variable_173_to_check;

// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_173[17:12] = value_check_98_to_variable_173;
assign enable_check_to_variable_173[2] = enable_check_98_to_variable_173;
// 将变量节点173的输出与校验节点98的输入相连
assign value_variable_173_to_check_98 = value_variable_173_to_check[17:12];
assign enable_variable_173_to_check_98 = enable_variable_173_to_check;


// 变量节点174的接口
wire [17:0] value_check_to_variable_174;
wire [2:0] enable_check_to_variable_174;
wire [5:0] value_variable_174_to_decision;
wire [17:0] value_variable_174_to_check;

wire enable_variable_174_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_174[5:0] = value_check_2_to_variable_174;
assign enable_check_to_variable_174[0] = enable_check_2_to_variable_174;
// 将变量节点174的输出与校验节点2的输入相连
assign value_variable_174_to_check_2 = value_variable_174_to_check[5:0];
assign enable_variable_174_to_check_2 = enable_variable_174_to_check;

// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_174[11:6] = value_check_53_to_variable_174;
assign enable_check_to_variable_174[1] = enable_check_53_to_variable_174;
// 将变量节点174的输出与校验节点53的输入相连
assign value_variable_174_to_check_53 = value_variable_174_to_check[11:6];
assign enable_variable_174_to_check_53 = enable_variable_174_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_174[17:12] = value_check_88_to_variable_174;
assign enable_check_to_variable_174[2] = enable_check_88_to_variable_174;
// 将变量节点174的输出与校验节点88的输入相连
assign value_variable_174_to_check_88 = value_variable_174_to_check[17:12];
assign enable_variable_174_to_check_88 = enable_variable_174_to_check;


// 变量节点175的接口
wire [17:0] value_check_to_variable_175;
wire [2:0] enable_check_to_variable_175;
wire [5:0] value_variable_175_to_decision;
wire [17:0] value_variable_175_to_check;

wire enable_variable_175_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_175[5:0] = value_check_3_to_variable_175;
assign enable_check_to_variable_175[0] = enable_check_3_to_variable_175;
// 将变量节点175的输出与校验节点3的输入相连
assign value_variable_175_to_check_3 = value_variable_175_to_check[5:0];
assign enable_variable_175_to_check_3 = enable_variable_175_to_check;

// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_175[11:6] = value_check_62_to_variable_175;
assign enable_check_to_variable_175[1] = enable_check_62_to_variable_175;
// 将变量节点175的输出与校验节点62的输入相连
assign value_variable_175_to_check_62 = value_variable_175_to_check[11:6];
assign enable_variable_175_to_check_62 = enable_variable_175_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_175[17:12] = value_check_126_to_variable_175;
assign enable_check_to_variable_175[2] = enable_check_126_to_variable_175;
// 将变量节点175的输出与校验节点126的输入相连
assign value_variable_175_to_check_126 = value_variable_175_to_check[17:12];
assign enable_variable_175_to_check_126 = enable_variable_175_to_check;


// 变量节点176的接口
wire [17:0] value_check_to_variable_176;
wire [2:0] enable_check_to_variable_176;
wire [5:0] value_variable_176_to_decision;
wire [17:0] value_variable_176_to_check;

wire enable_variable_176_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_176[5:0] = value_check_4_to_variable_176;
assign enable_check_to_variable_176[0] = enable_check_4_to_variable_176;
// 将变量节点176的输出与校验节点4的输入相连
assign value_variable_176_to_check_4 = value_variable_176_to_check[5:0];
assign enable_variable_176_to_check_4 = enable_variable_176_to_check;

// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_176[11:6] = value_check_43_to_variable_176;
assign enable_check_to_variable_176[1] = enable_check_43_to_variable_176;
// 将变量节点176的输出与校验节点43的输入相连
assign value_variable_176_to_check_43 = value_variable_176_to_check[11:6];
assign enable_variable_176_to_check_43 = enable_variable_176_to_check;

// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_176[17:12] = value_check_82_to_variable_176;
assign enable_check_to_variable_176[2] = enable_check_82_to_variable_176;
// 将变量节点176的输出与校验节点82的输入相连
assign value_variable_176_to_check_82 = value_variable_176_to_check[17:12];
assign enable_variable_176_to_check_82 = enable_variable_176_to_check;


// 变量节点177的接口
wire [17:0] value_check_to_variable_177;
wire [2:0] enable_check_to_variable_177;
wire [5:0] value_variable_177_to_decision;
wire [17:0] value_variable_177_to_check;

wire enable_variable_177_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_177[5:0] = value_check_5_to_variable_177;
assign enable_check_to_variable_177[0] = enable_check_5_to_variable_177;
// 将变量节点177的输出与校验节点5的输入相连
assign value_variable_177_to_check_5 = value_variable_177_to_check[5:0];
assign enable_variable_177_to_check_5 = enable_variable_177_to_check;

// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_177[11:6] = value_check_55_to_variable_177;
assign enable_check_to_variable_177[1] = enable_check_55_to_variable_177;
// 将变量节点177的输出与校验节点55的输入相连
assign value_variable_177_to_check_55 = value_variable_177_to_check[11:6];
assign enable_variable_177_to_check_55 = enable_variable_177_to_check;

// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_177[17:12] = value_check_69_to_variable_177;
assign enable_check_to_variable_177[2] = enable_check_69_to_variable_177;
// 将变量节点177的输出与校验节点69的输入相连
assign value_variable_177_to_check_69 = value_variable_177_to_check[17:12];
assign enable_variable_177_to_check_69 = enable_variable_177_to_check;


// 变量节点178的接口
wire [17:0] value_check_to_variable_178;
wire [2:0] enable_check_to_variable_178;
wire [5:0] value_variable_178_to_decision;
wire [17:0] value_variable_178_to_check;

wire enable_variable_178_to_check;
// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_178[5:0] = value_check_6_to_variable_178;
assign enable_check_to_variable_178[0] = enable_check_6_to_variable_178;
// 将变量节点178的输出与校验节点6的输入相连
assign value_variable_178_to_check_6 = value_variable_178_to_check[5:0];
assign enable_variable_178_to_check_6 = enable_variable_178_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_178[11:6] = value_check_96_to_variable_178;
assign enable_check_to_variable_178[1] = enable_check_96_to_variable_178;
// 将变量节点178的输出与校验节点96的输入相连
assign value_variable_178_to_check_96 = value_variable_178_to_check[11:6];
assign enable_variable_178_to_check_96 = enable_variable_178_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_178[17:12] = value_check_112_to_variable_178;
assign enable_check_to_variable_178[2] = enable_check_112_to_variable_178;
// 将变量节点178的输出与校验节点112的输入相连
assign value_variable_178_to_check_112 = value_variable_178_to_check[17:12];
assign enable_variable_178_to_check_112 = enable_variable_178_to_check;


// 变量节点179的接口
wire [17:0] value_check_to_variable_179;
wire [2:0] enable_check_to_variable_179;
wire [5:0] value_variable_179_to_decision;
wire [17:0] value_variable_179_to_check;

wire enable_variable_179_to_check;
// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_179[5:0] = value_check_7_to_variable_179;
assign enable_check_to_variable_179[0] = enable_check_7_to_variable_179;
// 将变量节点179的输出与校验节点7的输入相连
assign value_variable_179_to_check_7 = value_variable_179_to_check[5:0];
assign enable_variable_179_to_check_7 = enable_variable_179_to_check;

// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_179[11:6] = value_check_9_to_variable_179;
assign enable_check_to_variable_179[1] = enable_check_9_to_variable_179;
// 将变量节点179的输出与校验节点9的输入相连
assign value_variable_179_to_check_9 = value_variable_179_to_check[11:6];
assign enable_variable_179_to_check_9 = enable_variable_179_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_179[17:12] = value_check_117_to_variable_179;
assign enable_check_to_variable_179[2] = enable_check_117_to_variable_179;
// 将变量节点179的输出与校验节点117的输入相连
assign value_variable_179_to_check_117 = value_variable_179_to_check[17:12];
assign enable_variable_179_to_check_117 = enable_variable_179_to_check;


// 变量节点180的接口
wire [17:0] value_check_to_variable_180;
wire [2:0] enable_check_to_variable_180;
wire [5:0] value_variable_180_to_decision;
wire [17:0] value_variable_180_to_check;

wire enable_variable_180_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_180[5:0] = value_check_8_to_variable_180;
assign enable_check_to_variable_180[0] = enable_check_8_to_variable_180;
// 将变量节点180的输出与校验节点8的输入相连
assign value_variable_180_to_check_8 = value_variable_180_to_check[5:0];
assign enable_variable_180_to_check_8 = enable_variable_180_to_check;

// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_180[11:6] = value_check_29_to_variable_180;
assign enable_check_to_variable_180[1] = enable_check_29_to_variable_180;
// 将变量节点180的输出与校验节点29的输入相连
assign value_variable_180_to_check_29 = value_variable_180_to_check[11:6];
assign enable_variable_180_to_check_29 = enable_variable_180_to_check;

// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_180[17:12] = value_check_67_to_variable_180;
assign enable_check_to_variable_180[2] = enable_check_67_to_variable_180;
// 将变量节点180的输出与校验节点67的输入相连
assign value_variable_180_to_check_67 = value_variable_180_to_check[17:12];
assign enable_variable_180_to_check_67 = enable_variable_180_to_check;


// 变量节点181的接口
wire [17:0] value_check_to_variable_181;
wire [2:0] enable_check_to_variable_181;
wire [5:0] value_variable_181_to_decision;
wire [17:0] value_variable_181_to_check;

wire enable_variable_181_to_check;
// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_181[5:0] = value_check_10_to_variable_181;
assign enable_check_to_variable_181[0] = enable_check_10_to_variable_181;
// 将变量节点181的输出与校验节点10的输入相连
assign value_variable_181_to_check_10 = value_variable_181_to_check[5:0];
assign enable_variable_181_to_check_10 = enable_variable_181_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_181[11:6] = value_check_34_to_variable_181;
assign enable_check_to_variable_181[1] = enable_check_34_to_variable_181;
// 将变量节点181的输出与校验节点34的输入相连
assign value_variable_181_to_check_34 = value_variable_181_to_check[11:6];
assign enable_variable_181_to_check_34 = enable_variable_181_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_181[17:12] = value_check_101_to_variable_181;
assign enable_check_to_variable_181[2] = enable_check_101_to_variable_181;
// 将变量节点181的输出与校验节点101的输入相连
assign value_variable_181_to_check_101 = value_variable_181_to_check[17:12];
assign enable_variable_181_to_check_101 = enable_variable_181_to_check;


// 变量节点182的接口
wire [17:0] value_check_to_variable_182;
wire [2:0] enable_check_to_variable_182;
wire [5:0] value_variable_182_to_decision;
wire [17:0] value_variable_182_to_check;

wire enable_variable_182_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_182[5:0] = value_check_11_to_variable_182;
assign enable_check_to_variable_182[0] = enable_check_11_to_variable_182;
// 将变量节点182的输出与校验节点11的输入相连
assign value_variable_182_to_check_11 = value_variable_182_to_check[5:0];
assign enable_variable_182_to_check_11 = enable_variable_182_to_check;

// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_182[11:6] = value_check_24_to_variable_182;
assign enable_check_to_variable_182[1] = enable_check_24_to_variable_182;
// 将变量节点182的输出与校验节点24的输入相连
assign value_variable_182_to_check_24 = value_variable_182_to_check[11:6];
assign enable_variable_182_to_check_24 = enable_variable_182_to_check;

// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_182[17:12] = value_check_52_to_variable_182;
assign enable_check_to_variable_182[2] = enable_check_52_to_variable_182;
// 将变量节点182的输出与校验节点52的输入相连
assign value_variable_182_to_check_52 = value_variable_182_to_check[17:12];
assign enable_variable_182_to_check_52 = enable_variable_182_to_check;


// 变量节点183的接口
wire [17:0] value_check_to_variable_183;
wire [2:0] enable_check_to_variable_183;
wire [5:0] value_variable_183_to_decision;
wire [17:0] value_variable_183_to_check;

wire enable_variable_183_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_183[5:0] = value_check_12_to_variable_183;
assign enable_check_to_variable_183[0] = enable_check_12_to_variable_183;
// 将变量节点183的输出与校验节点12的输入相连
assign value_variable_183_to_check_12 = value_variable_183_to_check[5:0];
assign enable_variable_183_to_check_12 = enable_variable_183_to_check;

// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_183[11:6] = value_check_49_to_variable_183;
assign enable_check_to_variable_183[1] = enable_check_49_to_variable_183;
// 将变量节点183的输出与校验节点49的输入相连
assign value_variable_183_to_check_49 = value_variable_183_to_check[11:6];
assign enable_variable_183_to_check_49 = enable_variable_183_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_183[17:12] = value_check_85_to_variable_183;
assign enable_check_to_variable_183[2] = enable_check_85_to_variable_183;
// 将变量节点183的输出与校验节点85的输入相连
assign value_variable_183_to_check_85 = value_variable_183_to_check[17:12];
assign enable_variable_183_to_check_85 = enable_variable_183_to_check;


// 变量节点184的接口
wire [17:0] value_check_to_variable_184;
wire [2:0] enable_check_to_variable_184;
wire [5:0] value_variable_184_to_decision;
wire [17:0] value_variable_184_to_check;

wire enable_variable_184_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_184[5:0] = value_check_13_to_variable_184;
assign enable_check_to_variable_184[0] = enable_check_13_to_variable_184;
// 将变量节点184的输出与校验节点13的输入相连
assign value_variable_184_to_check_13 = value_variable_184_to_check[5:0];
assign enable_variable_184_to_check_13 = enable_variable_184_to_check;

// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_184[11:6] = value_check_16_to_variable_184;
assign enable_check_to_variable_184[1] = enable_check_16_to_variable_184;
// 将变量节点184的输出与校验节点16的输入相连
assign value_variable_184_to_check_16 = value_variable_184_to_check[11:6];
assign enable_variable_184_to_check_16 = enable_variable_184_to_check;

// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_184[17:12] = value_check_109_to_variable_184;
assign enable_check_to_variable_184[2] = enable_check_109_to_variable_184;
// 将变量节点184的输出与校验节点109的输入相连
assign value_variable_184_to_check_109 = value_variable_184_to_check[17:12];
assign enable_variable_184_to_check_109 = enable_variable_184_to_check;


// 变量节点185的接口
wire [17:0] value_check_to_variable_185;
wire [2:0] enable_check_to_variable_185;
wire [5:0] value_variable_185_to_decision;
wire [17:0] value_variable_185_to_check;

wire enable_variable_185_to_check;
// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_185[5:0] = value_check_14_to_variable_185;
assign enable_check_to_variable_185[0] = enable_check_14_to_variable_185;
// 将变量节点185的输出与校验节点14的输入相连
assign value_variable_185_to_check_14 = value_variable_185_to_check[5:0];
assign enable_variable_185_to_check_14 = enable_variable_185_to_check;

// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_185[11:6] = value_check_48_to_variable_185;
assign enable_check_to_variable_185[1] = enable_check_48_to_variable_185;
// 将变量节点185的输出与校验节点48的输入相连
assign value_variable_185_to_check_48 = value_variable_185_to_check[11:6];
assign enable_variable_185_to_check_48 = enable_variable_185_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_185[17:12] = value_check_127_to_variable_185;
assign enable_check_to_variable_185[2] = enable_check_127_to_variable_185;
// 将变量节点185的输出与校验节点127的输入相连
assign value_variable_185_to_check_127 = value_variable_185_to_check[17:12];
assign enable_variable_185_to_check_127 = enable_variable_185_to_check;


// 变量节点186的接口
wire [17:0] value_check_to_variable_186;
wire [2:0] enable_check_to_variable_186;
wire [5:0] value_variable_186_to_decision;
wire [17:0] value_variable_186_to_check;

wire enable_variable_186_to_check;
// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_186[5:0] = value_check_15_to_variable_186;
assign enable_check_to_variable_186[0] = enable_check_15_to_variable_186;
// 将变量节点186的输出与校验节点15的输入相连
assign value_variable_186_to_check_15 = value_variable_186_to_check[5:0];
assign enable_variable_186_to_check_15 = enable_variable_186_to_check;

// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_186[11:6] = value_check_19_to_variable_186;
assign enable_check_to_variable_186[1] = enable_check_19_to_variable_186;
// 将变量节点186的输出与校验节点19的输入相连
assign value_variable_186_to_check_19 = value_variable_186_to_check[11:6];
assign enable_variable_186_to_check_19 = enable_variable_186_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_186[17:12] = value_check_78_to_variable_186;
assign enable_check_to_variable_186[2] = enable_check_78_to_variable_186;
// 将变量节点186的输出与校验节点78的输入相连
assign value_variable_186_to_check_78 = value_variable_186_to_check[17:12];
assign enable_variable_186_to_check_78 = enable_variable_186_to_check;


// 变量节点187的接口
wire [17:0] value_check_to_variable_187;
wire [2:0] enable_check_to_variable_187;
wire [5:0] value_variable_187_to_decision;
wire [17:0] value_variable_187_to_check;

wire enable_variable_187_to_check;
// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_187[5:0] = value_check_17_to_variable_187;
assign enable_check_to_variable_187[0] = enable_check_17_to_variable_187;
// 将变量节点187的输出与校验节点17的输入相连
assign value_variable_187_to_check_17 = value_variable_187_to_check[5:0];
assign enable_variable_187_to_check_17 = enable_variable_187_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_187[11:6] = value_check_111_to_variable_187;
assign enable_check_to_variable_187[1] = enable_check_111_to_variable_187;
// 将变量节点187的输出与校验节点111的输入相连
assign value_variable_187_to_check_111 = value_variable_187_to_check[11:6];
assign enable_variable_187_to_check_111 = enable_variable_187_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_187[17:12] = value_check_120_to_variable_187;
assign enable_check_to_variable_187[2] = enable_check_120_to_variable_187;
// 将变量节点187的输出与校验节点120的输入相连
assign value_variable_187_to_check_120 = value_variable_187_to_check[17:12];
assign enable_variable_187_to_check_120 = enable_variable_187_to_check;


// 变量节点188的接口
wire [17:0] value_check_to_variable_188;
wire [2:0] enable_check_to_variable_188;
wire [5:0] value_variable_188_to_decision;
wire [17:0] value_variable_188_to_check;

wire enable_variable_188_to_check;
// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_188[5:0] = value_check_18_to_variable_188;
assign enable_check_to_variable_188[0] = enable_check_18_to_variable_188;
// 将变量节点188的输出与校验节点18的输入相连
assign value_variable_188_to_check_18 = value_variable_188_to_check[5:0];
assign enable_variable_188_to_check_18 = enable_variable_188_to_check;

// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_188[11:6] = value_check_21_to_variable_188;
assign enable_check_to_variable_188[1] = enable_check_21_to_variable_188;
// 将变量节点188的输出与校验节点21的输入相连
assign value_variable_188_to_check_21 = value_variable_188_to_check[11:6];
assign enable_variable_188_to_check_21 = enable_variable_188_to_check;

// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_188[17:12] = value_check_74_to_variable_188;
assign enable_check_to_variable_188[2] = enable_check_74_to_variable_188;
// 将变量节点188的输出与校验节点74的输入相连
assign value_variable_188_to_check_74 = value_variable_188_to_check[17:12];
assign enable_variable_188_to_check_74 = enable_variable_188_to_check;


// 变量节点189的接口
wire [17:0] value_check_to_variable_189;
wire [2:0] enable_check_to_variable_189;
wire [5:0] value_variable_189_to_decision;
wire [17:0] value_variable_189_to_check;

wire enable_variable_189_to_check;
// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_189[5:0] = value_check_22_to_variable_189;
assign enable_check_to_variable_189[0] = enable_check_22_to_variable_189;
// 将变量节点189的输出与校验节点22的输入相连
assign value_variable_189_to_check_22 = value_variable_189_to_check[5:0];
assign enable_variable_189_to_check_22 = enable_variable_189_to_check;

// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_189[11:6] = value_check_33_to_variable_189;
assign enable_check_to_variable_189[1] = enable_check_33_to_variable_189;
// 将变量节点189的输出与校验节点33的输入相连
assign value_variable_189_to_check_33 = value_variable_189_to_check[11:6];
assign enable_variable_189_to_check_33 = enable_variable_189_to_check;

// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_189[17:12] = value_check_37_to_variable_189;
assign enable_check_to_variable_189[2] = enable_check_37_to_variable_189;
// 将变量节点189的输出与校验节点37的输入相连
assign value_variable_189_to_check_37 = value_variable_189_to_check[17:12];
assign enable_variable_189_to_check_37 = enable_variable_189_to_check;


// 变量节点190的接口
wire [17:0] value_check_to_variable_190;
wire [2:0] enable_check_to_variable_190;
wire [5:0] value_variable_190_to_decision;
wire [17:0] value_variable_190_to_check;

wire enable_variable_190_to_check;
// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_190[5:0] = value_check_23_to_variable_190;
assign enable_check_to_variable_190[0] = enable_check_23_to_variable_190;
// 将变量节点190的输出与校验节点23的输入相连
assign value_variable_190_to_check_23 = value_variable_190_to_check[5:0];
assign enable_variable_190_to_check_23 = enable_variable_190_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_190[11:6] = value_check_91_to_variable_190;
assign enable_check_to_variable_190[1] = enable_check_91_to_variable_190;
// 将变量节点190的输出与校验节点91的输入相连
assign value_variable_190_to_check_91 = value_variable_190_to_check[11:6];
assign enable_variable_190_to_check_91 = enable_variable_190_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_190[17:12] = value_check_119_to_variable_190;
assign enable_check_to_variable_190[2] = enable_check_119_to_variable_190;
// 将变量节点190的输出与校验节点119的输入相连
assign value_variable_190_to_check_119 = value_variable_190_to_check[17:12];
assign enable_variable_190_to_check_119 = enable_variable_190_to_check;


// 变量节点191的接口
wire [17:0] value_check_to_variable_191;
wire [2:0] enable_check_to_variable_191;
wire [5:0] value_variable_191_to_decision;
wire [17:0] value_variable_191_to_check;

wire enable_variable_191_to_check;
// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_191[5:0] = value_check_25_to_variable_191;
assign enable_check_to_variable_191[0] = enable_check_25_to_variable_191;
// 将变量节点191的输出与校验节点25的输入相连
assign value_variable_191_to_check_25 = value_variable_191_to_check[5:0];
assign enable_variable_191_to_check_25 = enable_variable_191_to_check;

// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_191[11:6] = value_check_71_to_variable_191;
assign enable_check_to_variable_191[1] = enable_check_71_to_variable_191;
// 将变量节点191的输出与校验节点71的输入相连
assign value_variable_191_to_check_71 = value_variable_191_to_check[11:6];
assign enable_variable_191_to_check_71 = enable_variable_191_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_191[17:12] = value_check_122_to_variable_191;
assign enable_check_to_variable_191[2] = enable_check_122_to_variable_191;
// 将变量节点191的输出与校验节点122的输入相连
assign value_variable_191_to_check_122 = value_variable_191_to_check[17:12];
assign enable_variable_191_to_check_122 = enable_variable_191_to_check;


// 变量节点192的接口
wire [17:0] value_check_to_variable_192;
wire [2:0] enable_check_to_variable_192;
wire [5:0] value_variable_192_to_decision;
wire [17:0] value_variable_192_to_check;

wire enable_variable_192_to_check;
// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_192[5:0] = value_check_26_to_variable_192;
assign enable_check_to_variable_192[0] = enable_check_26_to_variable_192;
// 将变量节点192的输出与校验节点26的输入相连
assign value_variable_192_to_check_26 = value_variable_192_to_check[5:0];
assign enable_variable_192_to_check_26 = enable_variable_192_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_192[11:6] = value_check_94_to_variable_192;
assign enable_check_to_variable_192[1] = enable_check_94_to_variable_192;
// 将变量节点192的输出与校验节点94的输入相连
assign value_variable_192_to_check_94 = value_variable_192_to_check[11:6];
assign enable_variable_192_to_check_94 = enable_variable_192_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_192[17:12] = value_check_103_to_variable_192;
assign enable_check_to_variable_192[2] = enable_check_103_to_variable_192;
// 将变量节点192的输出与校验节点103的输入相连
assign value_variable_192_to_check_103 = value_variable_192_to_check[17:12];
assign enable_variable_192_to_check_103 = enable_variable_192_to_check;


// 变量节点193的接口
wire [17:0] value_check_to_variable_193;
wire [2:0] enable_check_to_variable_193;
wire [5:0] value_variable_193_to_decision;
wire [17:0] value_variable_193_to_check;

wire enable_variable_193_to_check;
// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_193[5:0] = value_check_27_to_variable_193;
assign enable_check_to_variable_193[0] = enable_check_27_to_variable_193;
// 将变量节点193的输出与校验节点27的输入相连
assign value_variable_193_to_check_27 = value_variable_193_to_check[5:0];
assign enable_variable_193_to_check_27 = enable_variable_193_to_check;

// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_193[11:6] = value_check_54_to_variable_193;
assign enable_check_to_variable_193[1] = enable_check_54_to_variable_193;
// 将变量节点193的输出与校验节点54的输入相连
assign value_variable_193_to_check_54 = value_variable_193_to_check[11:6];
assign enable_variable_193_to_check_54 = enable_variable_193_to_check;

// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_193[17:12] = value_check_59_to_variable_193;
assign enable_check_to_variable_193[2] = enable_check_59_to_variable_193;
// 将变量节点193的输出与校验节点59的输入相连
assign value_variable_193_to_check_59 = value_variable_193_to_check[17:12];
assign enable_variable_193_to_check_59 = enable_variable_193_to_check;


// 变量节点194的接口
wire [17:0] value_check_to_variable_194;
wire [2:0] enable_check_to_variable_194;
wire [5:0] value_variable_194_to_decision;
wire [17:0] value_variable_194_to_check;

wire enable_variable_194_to_check;
// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_194[5:0] = value_check_28_to_variable_194;
assign enable_check_to_variable_194[0] = enable_check_28_to_variable_194;
// 将变量节点194的输出与校验节点28的输入相连
assign value_variable_194_to_check_28 = value_variable_194_to_check[5:0];
assign enable_variable_194_to_check_28 = enable_variable_194_to_check;

// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_194[11:6] = value_check_76_to_variable_194;
assign enable_check_to_variable_194[1] = enable_check_76_to_variable_194;
// 将变量节点194的输出与校验节点76的输入相连
assign value_variable_194_to_check_76 = value_variable_194_to_check[11:6];
assign enable_variable_194_to_check_76 = enable_variable_194_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_194[17:12] = value_check_115_to_variable_194;
assign enable_check_to_variable_194[2] = enable_check_115_to_variable_194;
// 将变量节点194的输出与校验节点115的输入相连
assign value_variable_194_to_check_115 = value_variable_194_to_check[17:12];
assign enable_variable_194_to_check_115 = enable_variable_194_to_check;


// 变量节点195的接口
wire [17:0] value_check_to_variable_195;
wire [2:0] enable_check_to_variable_195;
wire [5:0] value_variable_195_to_decision;
wire [17:0] value_variable_195_to_check;

wire enable_variable_195_to_check;
// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_195[5:0] = value_check_30_to_variable_195;
assign enable_check_to_variable_195[0] = enable_check_30_to_variable_195;
// 将变量节点195的输出与校验节点30的输入相连
assign value_variable_195_to_check_30 = value_variable_195_to_check[5:0];
assign enable_variable_195_to_check_30 = enable_variable_195_to_check;

// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_195[11:6] = value_check_31_to_variable_195;
assign enable_check_to_variable_195[1] = enable_check_31_to_variable_195;
// 将变量节点195的输出与校验节点31的输入相连
assign value_variable_195_to_check_31 = value_variable_195_to_check[11:6];
assign enable_variable_195_to_check_31 = enable_variable_195_to_check;

// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_195[17:12] = value_check_45_to_variable_195;
assign enable_check_to_variable_195[2] = enable_check_45_to_variable_195;
// 将变量节点195的输出与校验节点45的输入相连
assign value_variable_195_to_check_45 = value_variable_195_to_check[17:12];
assign enable_variable_195_to_check_45 = enable_variable_195_to_check;


// 变量节点196的接口
wire [17:0] value_check_to_variable_196;
wire [2:0] enable_check_to_variable_196;
wire [5:0] value_variable_196_to_decision;
wire [17:0] value_variable_196_to_check;

wire enable_variable_196_to_check;
// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_196[5:0] = value_check_32_to_variable_196;
assign enable_check_to_variable_196[0] = enable_check_32_to_variable_196;
// 将变量节点196的输出与校验节点32的输入相连
assign value_variable_196_to_check_32 = value_variable_196_to_check[5:0];
assign enable_variable_196_to_check_32 = enable_variable_196_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_196[11:6] = value_check_89_to_variable_196;
assign enable_check_to_variable_196[1] = enable_check_89_to_variable_196;
// 将变量节点196的输出与校验节点89的输入相连
assign value_variable_196_to_check_89 = value_variable_196_to_check[11:6];
assign enable_variable_196_to_check_89 = enable_variable_196_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_196[17:12] = value_check_102_to_variable_196;
assign enable_check_to_variable_196[2] = enable_check_102_to_variable_196;
// 将变量节点196的输出与校验节点102的输入相连
assign value_variable_196_to_check_102 = value_variable_196_to_check[17:12];
assign enable_variable_196_to_check_102 = enable_variable_196_to_check;


// 变量节点197的接口
wire [17:0] value_check_to_variable_197;
wire [2:0] enable_check_to_variable_197;
wire [5:0] value_variable_197_to_decision;
wire [17:0] value_variable_197_to_check;

wire enable_variable_197_to_check;
// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_197[5:0] = value_check_35_to_variable_197;
assign enable_check_to_variable_197[0] = enable_check_35_to_variable_197;
// 将变量节点197的输出与校验节点35的输入相连
assign value_variable_197_to_check_35 = value_variable_197_to_check[5:0];
assign enable_variable_197_to_check_35 = enable_variable_197_to_check;

// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_197[11:6] = value_check_65_to_variable_197;
assign enable_check_to_variable_197[1] = enable_check_65_to_variable_197;
// 将变量节点197的输出与校验节点65的输入相连
assign value_variable_197_to_check_65 = value_variable_197_to_check[11:6];
assign enable_variable_197_to_check_65 = enable_variable_197_to_check;

// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_197[17:12] = value_check_70_to_variable_197;
assign enable_check_to_variable_197[2] = enable_check_70_to_variable_197;
// 将变量节点197的输出与校验节点70的输入相连
assign value_variable_197_to_check_70 = value_variable_197_to_check[17:12];
assign enable_variable_197_to_check_70 = enable_variable_197_to_check;


// 变量节点198的接口
wire [17:0] value_check_to_variable_198;
wire [2:0] enable_check_to_variable_198;
wire [5:0] value_variable_198_to_decision;
wire [17:0] value_variable_198_to_check;

wire enable_variable_198_to_check;
// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_198[5:0] = value_check_36_to_variable_198;
assign enable_check_to_variable_198[0] = enable_check_36_to_variable_198;
// 将变量节点198的输出与校验节点36的输入相连
assign value_variable_198_to_check_36 = value_variable_198_to_check[5:0];
assign enable_variable_198_to_check_36 = enable_variable_198_to_check;

// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_198[11:6] = value_check_47_to_variable_198;
assign enable_check_to_variable_198[1] = enable_check_47_to_variable_198;
// 将变量节点198的输出与校验节点47的输入相连
assign value_variable_198_to_check_47 = value_variable_198_to_check[11:6];
assign enable_variable_198_to_check_47 = enable_variable_198_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_198[17:12] = value_check_116_to_variable_198;
assign enable_check_to_variable_198[2] = enable_check_116_to_variable_198;
// 将变量节点198的输出与校验节点116的输入相连
assign value_variable_198_to_check_116 = value_variable_198_to_check[17:12];
assign enable_variable_198_to_check_116 = enable_variable_198_to_check;


// 变量节点199的接口
wire [17:0] value_check_to_variable_199;
wire [2:0] enable_check_to_variable_199;
wire [5:0] value_variable_199_to_decision;
wire [17:0] value_variable_199_to_check;

wire enable_variable_199_to_check;
// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_199[5:0] = value_check_39_to_variable_199;
assign enable_check_to_variable_199[0] = enable_check_39_to_variable_199;
// 将变量节点199的输出与校验节点39的输入相连
assign value_variable_199_to_check_39 = value_variable_199_to_check[5:0];
assign enable_variable_199_to_check_39 = enable_variable_199_to_check;

// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_199[11:6] = value_check_66_to_variable_199;
assign enable_check_to_variable_199[1] = enable_check_66_to_variable_199;
// 将变量节点199的输出与校验节点66的输入相连
assign value_variable_199_to_check_66 = value_variable_199_to_check[11:6];
assign enable_variable_199_to_check_66 = enable_variable_199_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_199[17:12] = value_check_93_to_variable_199;
assign enable_check_to_variable_199[2] = enable_check_93_to_variable_199;
// 将变量节点199的输出与校验节点93的输入相连
assign value_variable_199_to_check_93 = value_variable_199_to_check[17:12];
assign enable_variable_199_to_check_93 = enable_variable_199_to_check;


// 变量节点200的接口
wire [17:0] value_check_to_variable_200;
wire [2:0] enable_check_to_variable_200;
wire [5:0] value_variable_200_to_decision;
wire [17:0] value_variable_200_to_check;

wire enable_variable_200_to_check;
// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_200[5:0] = value_check_40_to_variable_200;
assign enable_check_to_variable_200[0] = enable_check_40_to_variable_200;
// 将变量节点200的输出与校验节点40的输入相连
assign value_variable_200_to_check_40 = value_variable_200_to_check[5:0];
assign enable_variable_200_to_check_40 = enable_variable_200_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_200[11:6] = value_check_75_to_variable_200;
assign enable_check_to_variable_200[1] = enable_check_75_to_variable_200;
// 将变量节点200的输出与校验节点75的输入相连
assign value_variable_200_to_check_75 = value_variable_200_to_check[11:6];
assign enable_variable_200_to_check_75 = enable_variable_200_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_200[17:12] = value_check_106_to_variable_200;
assign enable_check_to_variable_200[2] = enable_check_106_to_variable_200;
// 将变量节点200的输出与校验节点106的输入相连
assign value_variable_200_to_check_106 = value_variable_200_to_check[17:12];
assign enable_variable_200_to_check_106 = enable_variable_200_to_check;


// 变量节点201的接口
wire [17:0] value_check_to_variable_201;
wire [2:0] enable_check_to_variable_201;
wire [5:0] value_variable_201_to_decision;
wire [17:0] value_variable_201_to_check;

wire enable_variable_201_to_check;
// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_201[5:0] = value_check_41_to_variable_201;
assign enable_check_to_variable_201[0] = enable_check_41_to_variable_201;
// 将变量节点201的输出与校验节点41的输入相连
assign value_variable_201_to_check_41 = value_variable_201_to_check[5:0];
assign enable_variable_201_to_check_41 = enable_variable_201_to_check;

// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_201[11:6] = value_check_80_to_variable_201;
assign enable_check_to_variable_201[1] = enable_check_80_to_variable_201;
// 将变量节点201的输出与校验节点80的输入相连
assign value_variable_201_to_check_80 = value_variable_201_to_check[11:6];
assign enable_variable_201_to_check_80 = enable_variable_201_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_201[17:12] = value_check_81_to_variable_201;
assign enable_check_to_variable_201[2] = enable_check_81_to_variable_201;
// 将变量节点201的输出与校验节点81的输入相连
assign value_variable_201_to_check_81 = value_variable_201_to_check[17:12];
assign enable_variable_201_to_check_81 = enable_variable_201_to_check;


// 变量节点202的接口
wire [17:0] value_check_to_variable_202;
wire [2:0] enable_check_to_variable_202;
wire [5:0] value_variable_202_to_decision;
wire [17:0] value_variable_202_to_check;

wire enable_variable_202_to_check;
// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_202[5:0] = value_check_42_to_variable_202;
assign enable_check_to_variable_202[0] = enable_check_42_to_variable_202;
// 将变量节点202的输出与校验节点42的输入相连
assign value_variable_202_to_check_42 = value_variable_202_to_check[5:0];
assign enable_variable_202_to_check_42 = enable_variable_202_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_202[11:6] = value_check_61_to_variable_202;
assign enable_check_to_variable_202[1] = enable_check_61_to_variable_202;
// 将变量节点202的输出与校验节点61的输入相连
assign value_variable_202_to_check_61 = value_variable_202_to_check[11:6];
assign enable_variable_202_to_check_61 = enable_variable_202_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_202[17:12] = value_check_123_to_variable_202;
assign enable_check_to_variable_202[2] = enable_check_123_to_variable_202;
// 将变量节点202的输出与校验节点123的输入相连
assign value_variable_202_to_check_123 = value_variable_202_to_check[17:12];
assign enable_variable_202_to_check_123 = enable_variable_202_to_check;


// 变量节点203的接口
wire [17:0] value_check_to_variable_203;
wire [2:0] enable_check_to_variable_203;
wire [5:0] value_variable_203_to_decision;
wire [17:0] value_variable_203_to_check;

wire enable_variable_203_to_check;
// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_203[5:0] = value_check_44_to_variable_203;
assign enable_check_to_variable_203[0] = enable_check_44_to_variable_203;
// 将变量节点203的输出与校验节点44的输入相连
assign value_variable_203_to_check_44 = value_variable_203_to_check[5:0];
assign enable_variable_203_to_check_44 = enable_variable_203_to_check;

// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_203[11:6] = value_check_83_to_variable_203;
assign enable_check_to_variable_203[1] = enable_check_83_to_variable_203;
// 将变量节点203的输出与校验节点83的输入相连
assign value_variable_203_to_check_83 = value_variable_203_to_check[11:6];
assign enable_variable_203_to_check_83 = enable_variable_203_to_check;

// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_203[17:12] = value_check_100_to_variable_203;
assign enable_check_to_variable_203[2] = enable_check_100_to_variable_203;
// 将变量节点203的输出与校验节点100的输入相连
assign value_variable_203_to_check_100 = value_variable_203_to_check[17:12];
assign enable_variable_203_to_check_100 = enable_variable_203_to_check;


// 变量节点204的接口
wire [17:0] value_check_to_variable_204;
wire [2:0] enable_check_to_variable_204;
wire [5:0] value_variable_204_to_decision;
wire [17:0] value_variable_204_to_check;

wire enable_variable_204_to_check;
// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_204[5:0] = value_check_46_to_variable_204;
assign enable_check_to_variable_204[0] = enable_check_46_to_variable_204;
// 将变量节点204的输出与校验节点46的输入相连
assign value_variable_204_to_check_46 = value_variable_204_to_check[5:0];
assign enable_variable_204_to_check_46 = enable_variable_204_to_check;

// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_204[11:6] = value_check_58_to_variable_204;
assign enable_check_to_variable_204[1] = enable_check_58_to_variable_204;
// 将变量节点204的输出与校验节点58的输入相连
assign value_variable_204_to_check_58 = value_variable_204_to_check[11:6];
assign enable_variable_204_to_check_58 = enable_variable_204_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_204[17:12] = value_check_105_to_variable_204;
assign enable_check_to_variable_204[2] = enable_check_105_to_variable_204;
// 将变量节点204的输出与校验节点105的输入相连
assign value_variable_204_to_check_105 = value_variable_204_to_check[17:12];
assign enable_variable_204_to_check_105 = enable_variable_204_to_check;


// 变量节点205的接口
wire [17:0] value_check_to_variable_205;
wire [2:0] enable_check_to_variable_205;
wire [5:0] value_variable_205_to_decision;
wire [17:0] value_variable_205_to_check;

wire enable_variable_205_to_check;
// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_205[5:0] = value_check_51_to_variable_205;
assign enable_check_to_variable_205[0] = enable_check_51_to_variable_205;
// 将变量节点205的输出与校验节点51的输入相连
assign value_variable_205_to_check_51 = value_variable_205_to_check[5:0];
assign enable_variable_205_to_check_51 = enable_variable_205_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_205[11:6] = value_check_77_to_variable_205;
assign enable_check_to_variable_205[1] = enable_check_77_to_variable_205;
// 将变量节点205的输出与校验节点77的输入相连
assign value_variable_205_to_check_77 = value_variable_205_to_check[11:6];
assign enable_variable_205_to_check_77 = enable_variable_205_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_205[17:12] = value_check_104_to_variable_205;
assign enable_check_to_variable_205[2] = enable_check_104_to_variable_205;
// 将变量节点205的输出与校验节点104的输入相连
assign value_variable_205_to_check_104 = value_variable_205_to_check[17:12];
assign enable_variable_205_to_check_104 = enable_variable_205_to_check;


// 变量节点206的接口
wire [17:0] value_check_to_variable_206;
wire [2:0] enable_check_to_variable_206;
wire [5:0] value_variable_206_to_decision;
wire [17:0] value_variable_206_to_check;

wire enable_variable_206_to_check;
// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_206[5:0] = value_check_56_to_variable_206;
assign enable_check_to_variable_206[0] = enable_check_56_to_variable_206;
// 将变量节点206的输出与校验节点56的输入相连
assign value_variable_206_to_check_56 = value_variable_206_to_check[5:0];
assign enable_variable_206_to_check_56 = enable_variable_206_to_check;

// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_206[11:6] = value_check_72_to_variable_206;
assign enable_check_to_variable_206[1] = enable_check_72_to_variable_206;
// 将变量节点206的输出与校验节点72的输入相连
assign value_variable_206_to_check_72 = value_variable_206_to_check[11:6];
assign enable_variable_206_to_check_72 = enable_variable_206_to_check;

// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_206[17:12] = value_check_110_to_variable_206;
assign enable_check_to_variable_206[2] = enable_check_110_to_variable_206;
// 将变量节点206的输出与校验节点110的输入相连
assign value_variable_206_to_check_110 = value_variable_206_to_check[17:12];
assign enable_variable_206_to_check_110 = enable_variable_206_to_check;


// 变量节点207的接口
wire [17:0] value_check_to_variable_207;
wire [2:0] enable_check_to_variable_207;
wire [5:0] value_variable_207_to_decision;
wire [17:0] value_variable_207_to_check;

wire enable_variable_207_to_check;
// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_207[5:0] = value_check_63_to_variable_207;
assign enable_check_to_variable_207[0] = enable_check_63_to_variable_207;
// 将变量节点207的输出与校验节点63的输入相连
assign value_variable_207_to_check_63 = value_variable_207_to_check[5:0];
assign enable_variable_207_to_check_63 = enable_variable_207_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_207[11:6] = value_check_90_to_variable_207;
assign enable_check_to_variable_207[1] = enable_check_90_to_variable_207;
// 将变量节点207的输出与校验节点90的输入相连
assign value_variable_207_to_check_90 = value_variable_207_to_check[11:6];
assign enable_variable_207_to_check_90 = enable_variable_207_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_207[17:12] = value_check_92_to_variable_207;
assign enable_check_to_variable_207[2] = enable_check_92_to_variable_207;
// 将变量节点207的输出与校验节点92的输入相连
assign value_variable_207_to_check_92 = value_variable_207_to_check[17:12];
assign enable_variable_207_to_check_92 = enable_variable_207_to_check;


// 变量节点208的接口
wire [17:0] value_check_to_variable_208;
wire [2:0] enable_check_to_variable_208;
wire [5:0] value_variable_208_to_decision;
wire [17:0] value_variable_208_to_check;

wire enable_variable_208_to_check;
// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_208[5:0] = value_check_68_to_variable_208;
assign enable_check_to_variable_208[0] = enable_check_68_to_variable_208;
// 将变量节点208的输出与校验节点68的输入相连
assign value_variable_208_to_check_68 = value_variable_208_to_check[5:0];
assign enable_variable_208_to_check_68 = enable_variable_208_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_208[11:6] = value_check_87_to_variable_208;
assign enable_check_to_variable_208[1] = enable_check_87_to_variable_208;
// 将变量节点208的输出与校验节点87的输入相连
assign value_variable_208_to_check_87 = value_variable_208_to_check[11:6];
assign enable_variable_208_to_check_87 = enable_variable_208_to_check;

// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_208[17:12] = value_check_95_to_variable_208;
assign enable_check_to_variable_208[2] = enable_check_95_to_variable_208;
// 将变量节点208的输出与校验节点95的输入相连
assign value_variable_208_to_check_95 = value_variable_208_to_check[17:12];
assign enable_variable_208_to_check_95 = enable_variable_208_to_check;


// 变量节点209的接口
wire [17:0] value_check_to_variable_209;
wire [2:0] enable_check_to_variable_209;
wire [5:0] value_variable_209_to_decision;
wire [17:0] value_variable_209_to_check;

wire enable_variable_209_to_check;
// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_209[5:0] = value_check_73_to_variable_209;
assign enable_check_to_variable_209[0] = enable_check_73_to_variable_209;
// 将变量节点209的输出与校验节点73的输入相连
assign value_variable_209_to_check_73 = value_variable_209_to_check[5:0];
assign enable_variable_209_to_check_73 = enable_variable_209_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_209[11:6] = value_check_84_to_variable_209;
assign enable_check_to_variable_209[1] = enable_check_84_to_variable_209;
// 将变量节点209的输出与校验节点84的输入相连
assign value_variable_209_to_check_84 = value_variable_209_to_check[11:6];
assign enable_variable_209_to_check_84 = enable_variable_209_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_209[17:12] = value_check_121_to_variable_209;
assign enable_check_to_variable_209[2] = enable_check_121_to_variable_209;
// 将变量节点209的输出与校验节点121的输入相连
assign value_variable_209_to_check_121 = value_variable_209_to_check[17:12];
assign enable_variable_209_to_check_121 = enable_variable_209_to_check;


// 变量节点210的接口
wire [17:0] value_check_to_variable_210;
wire [2:0] enable_check_to_variable_210;
wire [5:0] value_variable_210_to_decision;
wire [17:0] value_variable_210_to_check;

wire enable_variable_210_to_check;
// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_210[5:0] = value_check_79_to_variable_210;
assign enable_check_to_variable_210[0] = enable_check_79_to_variable_210;
// 将变量节点210的输出与校验节点79的输入相连
assign value_variable_210_to_check_79 = value_variable_210_to_check[5:0];
assign enable_variable_210_to_check_79 = enable_variable_210_to_check;

// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_210[11:6] = value_check_86_to_variable_210;
assign enable_check_to_variable_210[1] = enable_check_86_to_variable_210;
// 将变量节点210的输出与校验节点86的输入相连
assign value_variable_210_to_check_86 = value_variable_210_to_check[11:6];
assign enable_variable_210_to_check_86 = enable_variable_210_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_210[17:12] = value_check_108_to_variable_210;
assign enable_check_to_variable_210[2] = enable_check_108_to_variable_210;
// 将变量节点210的输出与校验节点108的输入相连
assign value_variable_210_to_check_108 = value_variable_210_to_check[17:12];
assign enable_variable_210_to_check_108 = enable_variable_210_to_check;


// 变量节点211的接口
wire [17:0] value_check_to_variable_211;
wire [2:0] enable_check_to_variable_211;
wire [5:0] value_variable_211_to_decision;
wire [17:0] value_variable_211_to_check;

wire enable_variable_211_to_check;
// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_211[5:0] = value_check_97_to_variable_211;
assign enable_check_to_variable_211[0] = enable_check_97_to_variable_211;
// 将变量节点211的输出与校验节点97的输入相连
assign value_variable_211_to_check_97 = value_variable_211_to_check[5:0];
assign enable_variable_211_to_check_97 = enable_variable_211_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_211[11:6] = value_check_114_to_variable_211;
assign enable_check_to_variable_211[1] = enable_check_114_to_variable_211;
// 将变量节点211的输出与校验节点114的输入相连
assign value_variable_211_to_check_114 = value_variable_211_to_check[11:6];
assign enable_variable_211_to_check_114 = enable_variable_211_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_211[17:12] = value_check_124_to_variable_211;
assign enable_check_to_variable_211[2] = enable_check_124_to_variable_211;
// 将变量节点211的输出与校验节点124的输入相连
assign value_variable_211_to_check_124 = value_variable_211_to_check[17:12];
assign enable_variable_211_to_check_124 = enable_variable_211_to_check;


// 变量节点212的接口
wire [17:0] value_check_to_variable_212;
wire [2:0] enable_check_to_variable_212;
wire [5:0] value_variable_212_to_decision;
wire [17:0] value_variable_212_to_check;

wire enable_variable_212_to_check;
// 对校验节点69传递过来的数据进行整合
assign value_check_to_variable_212[5:0] = value_check_69_to_variable_212;
assign enable_check_to_variable_212[0] = enable_check_69_to_variable_212;
// 将变量节点212的输出与校验节点69的输入相连
assign value_variable_212_to_check_69 = value_variable_212_to_check[5:0];
assign enable_variable_212_to_check_69 = enable_variable_212_to_check;

// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_212[11:6] = value_check_99_to_variable_212;
assign enable_check_to_variable_212[1] = enable_check_99_to_variable_212;
// 将变量节点212的输出与校验节点99的输入相连
assign value_variable_212_to_check_99 = value_variable_212_to_check[11:6];
assign enable_variable_212_to_check_99 = enable_variable_212_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_212[17:12] = value_check_125_to_variable_212;
assign enable_check_to_variable_212[2] = enable_check_125_to_variable_212;
// 将变量节点212的输出与校验节点125的输入相连
assign value_variable_212_to_check_125 = value_variable_212_to_check[17:12];
assign enable_variable_212_to_check_125 = enable_variable_212_to_check;


// 变量节点213的接口
wire [17:0] value_check_to_variable_213;
wire [2:0] enable_check_to_variable_213;
wire [5:0] value_variable_213_to_decision;
wire [17:0] value_variable_213_to_check;

wire enable_variable_213_to_check;
// 对校验节点37传递过来的数据进行整合
assign value_check_to_variable_213[5:0] = value_check_37_to_variable_213;
assign enable_check_to_variable_213[0] = enable_check_37_to_variable_213;
// 将变量节点213的输出与校验节点37的输入相连
assign value_variable_213_to_check_37 = value_variable_213_to_check[5:0];
assign enable_variable_213_to_check_37 = enable_variable_213_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_213[11:6] = value_check_107_to_variable_213;
assign enable_check_to_variable_213[1] = enable_check_107_to_variable_213;
// 将变量节点213的输出与校验节点107的输入相连
assign value_variable_213_to_check_107 = value_variable_213_to_check[11:6];
assign enable_variable_213_to_check_107 = enable_variable_213_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_213[17:12] = value_check_113_to_variable_213;
assign enable_check_to_variable_213[2] = enable_check_113_to_variable_213;
// 将变量节点213的输出与校验节点113的输入相连
assign value_variable_213_to_check_113 = value_variable_213_to_check[17:12];
assign enable_variable_213_to_check_113 = enable_variable_213_to_check;


// 变量节点214的接口
wire [17:0] value_check_to_variable_214;
wire [2:0] enable_check_to_variable_214;
wire [5:0] value_variable_214_to_decision;
wire [17:0] value_variable_214_to_check;

wire enable_variable_214_to_check;
// 对校验节点0传递过来的数据进行整合
assign value_check_to_variable_214[5:0] = value_check_0_to_variable_214;
assign enable_check_to_variable_214[0] = enable_check_0_to_variable_214;
// 将变量节点214的输出与校验节点0的输入相连
assign value_variable_214_to_check_0 = value_variable_214_to_check[5:0];
assign enable_variable_214_to_check_0 = enable_variable_214_to_check;

// 对校验节点32传递过来的数据进行整合
assign value_check_to_variable_214[11:6] = value_check_32_to_variable_214;
assign enable_check_to_variable_214[1] = enable_check_32_to_variable_214;
// 将变量节点214的输出与校验节点32的输入相连
assign value_variable_214_to_check_32 = value_variable_214_to_check[11:6];
assign enable_variable_214_to_check_32 = enable_variable_214_to_check;

// 对校验节点117传递过来的数据进行整合
assign value_check_to_variable_214[17:12] = value_check_117_to_variable_214;
assign enable_check_to_variable_214[2] = enable_check_117_to_variable_214;
// 将变量节点214的输出与校验节点117的输入相连
assign value_variable_214_to_check_117 = value_variable_214_to_check[17:12];
assign enable_variable_214_to_check_117 = enable_variable_214_to_check;


// 变量节点215的接口
wire [17:0] value_check_to_variable_215;
wire [2:0] enable_check_to_variable_215;
wire [5:0] value_variable_215_to_decision;
wire [17:0] value_variable_215_to_check;

wire enable_variable_215_to_check;
// 对校验节点1传递过来的数据进行整合
assign value_check_to_variable_215[5:0] = value_check_1_to_variable_215;
assign enable_check_to_variable_215[0] = enable_check_1_to_variable_215;
// 将变量节点215的输出与校验节点1的输入相连
assign value_variable_215_to_check_1 = value_variable_215_to_check[5:0];
assign enable_variable_215_to_check_1 = enable_variable_215_to_check;

// 对校验节点99传递过来的数据进行整合
assign value_check_to_variable_215[11:6] = value_check_99_to_variable_215;
assign enable_check_to_variable_215[1] = enable_check_99_to_variable_215;
// 将变量节点215的输出与校验节点99的输入相连
assign value_variable_215_to_check_99 = value_variable_215_to_check[11:6];
assign enable_variable_215_to_check_99 = enable_variable_215_to_check;

// 对校验节点119传递过来的数据进行整合
assign value_check_to_variable_215[17:12] = value_check_119_to_variable_215;
assign enable_check_to_variable_215[2] = enable_check_119_to_variable_215;
// 将变量节点215的输出与校验节点119的输入相连
assign value_variable_215_to_check_119 = value_variable_215_to_check[17:12];
assign enable_variable_215_to_check_119 = enable_variable_215_to_check;


// 变量节点216的接口
wire [17:0] value_check_to_variable_216;
wire [2:0] enable_check_to_variable_216;
wire [5:0] value_variable_216_to_decision;
wire [17:0] value_variable_216_to_check;

wire enable_variable_216_to_check;
// 对校验节点2传递过来的数据进行整合
assign value_check_to_variable_216[5:0] = value_check_2_to_variable_216;
assign enable_check_to_variable_216[0] = enable_check_2_to_variable_216;
// 将变量节点216的输出与校验节点2的输入相连
assign value_variable_216_to_check_2 = value_variable_216_to_check[5:0];
assign enable_variable_216_to_check_2 = enable_variable_216_to_check;

// 对校验节点16传递过来的数据进行整合
assign value_check_to_variable_216[11:6] = value_check_16_to_variable_216;
assign enable_check_to_variable_216[1] = enable_check_16_to_variable_216;
// 将变量节点216的输出与校验节点16的输入相连
assign value_variable_216_to_check_16 = value_variable_216_to_check[11:6];
assign enable_variable_216_to_check_16 = enable_variable_216_to_check;

// 对校验节点73传递过来的数据进行整合
assign value_check_to_variable_216[17:12] = value_check_73_to_variable_216;
assign enable_check_to_variable_216[2] = enable_check_73_to_variable_216;
// 将变量节点216的输出与校验节点73的输入相连
assign value_variable_216_to_check_73 = value_variable_216_to_check[17:12];
assign enable_variable_216_to_check_73 = enable_variable_216_to_check;


// 变量节点217的接口
wire [17:0] value_check_to_variable_217;
wire [2:0] enable_check_to_variable_217;
wire [5:0] value_variable_217_to_decision;
wire [17:0] value_variable_217_to_check;

wire enable_variable_217_to_check;
// 对校验节点3传递过来的数据进行整合
assign value_check_to_variable_217[5:0] = value_check_3_to_variable_217;
assign enable_check_to_variable_217[0] = enable_check_3_to_variable_217;
// 将变量节点217的输出与校验节点3的输入相连
assign value_variable_217_to_check_3 = value_variable_217_to_check[5:0];
assign enable_variable_217_to_check_3 = enable_variable_217_to_check;

// 对校验节点15传递过来的数据进行整合
assign value_check_to_variable_217[11:6] = value_check_15_to_variable_217;
assign enable_check_to_variable_217[1] = enable_check_15_to_variable_217;
// 将变量节点217的输出与校验节点15的输入相连
assign value_variable_217_to_check_15 = value_variable_217_to_check[11:6];
assign enable_variable_217_to_check_15 = enable_variable_217_to_check;

// 对校验节点63传递过来的数据进行整合
assign value_check_to_variable_217[17:12] = value_check_63_to_variable_217;
assign enable_check_to_variable_217[2] = enable_check_63_to_variable_217;
// 将变量节点217的输出与校验节点63的输入相连
assign value_variable_217_to_check_63 = value_variable_217_to_check[17:12];
assign enable_variable_217_to_check_63 = enable_variable_217_to_check;


// 变量节点218的接口
wire [17:0] value_check_to_variable_218;
wire [2:0] enable_check_to_variable_218;
wire [5:0] value_variable_218_to_decision;
wire [17:0] value_variable_218_to_check;

wire enable_variable_218_to_check;
// 对校验节点4传递过来的数据进行整合
assign value_check_to_variable_218[5:0] = value_check_4_to_variable_218;
assign enable_check_to_variable_218[0] = enable_check_4_to_variable_218;
// 将变量节点218的输出与校验节点4的输入相连
assign value_variable_218_to_check_4 = value_variable_218_to_check[5:0];
assign enable_variable_218_to_check_4 = enable_variable_218_to_check;

// 对校验节点21传递过来的数据进行整合
assign value_check_to_variable_218[11:6] = value_check_21_to_variable_218;
assign enable_check_to_variable_218[1] = enable_check_21_to_variable_218;
// 将变量节点218的输出与校验节点21的输入相连
assign value_variable_218_to_check_21 = value_variable_218_to_check[11:6];
assign enable_variable_218_to_check_21 = enable_variable_218_to_check;

// 对校验节点78传递过来的数据进行整合
assign value_check_to_variable_218[17:12] = value_check_78_to_variable_218;
assign enable_check_to_variable_218[2] = enable_check_78_to_variable_218;
// 将变量节点218的输出与校验节点78的输入相连
assign value_variable_218_to_check_78 = value_variable_218_to_check[17:12];
assign enable_variable_218_to_check_78 = enable_variable_218_to_check;


// 变量节点219的接口
wire [17:0] value_check_to_variable_219;
wire [2:0] enable_check_to_variable_219;
wire [5:0] value_variable_219_to_decision;
wire [17:0] value_variable_219_to_check;

wire enable_variable_219_to_check;
// 对校验节点5传递过来的数据进行整合
assign value_check_to_variable_219[5:0] = value_check_5_to_variable_219;
assign enable_check_to_variable_219[0] = enable_check_5_to_variable_219;
// 将变量节点219的输出与校验节点5的输入相连
assign value_variable_219_to_check_5 = value_variable_219_to_check[5:0];
assign enable_variable_219_to_check_5 = enable_variable_219_to_check;

// 对校验节点43传递过来的数据进行整合
assign value_check_to_variable_219[11:6] = value_check_43_to_variable_219;
assign enable_check_to_variable_219[1] = enable_check_43_to_variable_219;
// 将变量节点219的输出与校验节点43的输入相连
assign value_variable_219_to_check_43 = value_variable_219_to_check[11:6];
assign enable_variable_219_to_check_43 = enable_variable_219_to_check;

// 对校验节点89传递过来的数据进行整合
assign value_check_to_variable_219[17:12] = value_check_89_to_variable_219;
assign enable_check_to_variable_219[2] = enable_check_89_to_variable_219;
// 将变量节点219的输出与校验节点89的输入相连
assign value_variable_219_to_check_89 = value_variable_219_to_check[17:12];
assign enable_variable_219_to_check_89 = enable_variable_219_to_check;


// 变量节点220的接口
wire [17:0] value_check_to_variable_220;
wire [2:0] enable_check_to_variable_220;
wire [5:0] value_variable_220_to_decision;
wire [17:0] value_variable_220_to_check;

wire enable_variable_220_to_check;
// 对校验节点6传递过来的数据进行整合
assign value_check_to_variable_220[5:0] = value_check_6_to_variable_220;
assign enable_check_to_variable_220[0] = enable_check_6_to_variable_220;
// 将变量节点220的输出与校验节点6的输入相连
assign value_variable_220_to_check_6 = value_variable_220_to_check[5:0];
assign enable_variable_220_to_check_6 = enable_variable_220_to_check;

// 对校验节点30传递过来的数据进行整合
assign value_check_to_variable_220[11:6] = value_check_30_to_variable_220;
assign enable_check_to_variable_220[1] = enable_check_30_to_variable_220;
// 将变量节点220的输出与校验节点30的输入相连
assign value_variable_220_to_check_30 = value_variable_220_to_check[11:6];
assign enable_variable_220_to_check_30 = enable_variable_220_to_check;

// 对校验节点83传递过来的数据进行整合
assign value_check_to_variable_220[17:12] = value_check_83_to_variable_220;
assign enable_check_to_variable_220[2] = enable_check_83_to_variable_220;
// 将变量节点220的输出与校验节点83的输入相连
assign value_variable_220_to_check_83 = value_variable_220_to_check[17:12];
assign enable_variable_220_to_check_83 = enable_variable_220_to_check;


// 变量节点221的接口
wire [17:0] value_check_to_variable_221;
wire [2:0] enable_check_to_variable_221;
wire [5:0] value_variable_221_to_decision;
wire [17:0] value_variable_221_to_check;

wire enable_variable_221_to_check;
// 对校验节点7传递过来的数据进行整合
assign value_check_to_variable_221[5:0] = value_check_7_to_variable_221;
assign enable_check_to_variable_221[0] = enable_check_7_to_variable_221;
// 将变量节点221的输出与校验节点7的输入相连
assign value_variable_221_to_check_7 = value_variable_221_to_check[5:0];
assign enable_variable_221_to_check_7 = enable_variable_221_to_check;

// 对校验节点38传递过来的数据进行整合
assign value_check_to_variable_221[11:6] = value_check_38_to_variable_221;
assign enable_check_to_variable_221[1] = enable_check_38_to_variable_221;
// 将变量节点221的输出与校验节点38的输入相连
assign value_variable_221_to_check_38 = value_variable_221_to_check[11:6];
assign enable_variable_221_to_check_38 = enable_variable_221_to_check;

// 对校验节点101传递过来的数据进行整合
assign value_check_to_variable_221[17:12] = value_check_101_to_variable_221;
assign enable_check_to_variable_221[2] = enable_check_101_to_variable_221;
// 将变量节点221的输出与校验节点101的输入相连
assign value_variable_221_to_check_101 = value_variable_221_to_check[17:12];
assign enable_variable_221_to_check_101 = enable_variable_221_to_check;


// 变量节点222的接口
wire [17:0] value_check_to_variable_222;
wire [2:0] enable_check_to_variable_222;
wire [5:0] value_variable_222_to_decision;
wire [17:0] value_variable_222_to_check;

wire enable_variable_222_to_check;
// 对校验节点8传递过来的数据进行整合
assign value_check_to_variable_222[5:0] = value_check_8_to_variable_222;
assign enable_check_to_variable_222[0] = enable_check_8_to_variable_222;
// 将变量节点222的输出与校验节点8的输入相连
assign value_variable_222_to_check_8 = value_variable_222_to_check[5:0];
assign enable_variable_222_to_check_8 = enable_variable_222_to_check;

// 对校验节点10传递过来的数据进行整合
assign value_check_to_variable_222[11:6] = value_check_10_to_variable_222;
assign enable_check_to_variable_222[1] = enable_check_10_to_variable_222;
// 将变量节点222的输出与校验节点10的输入相连
assign value_variable_222_to_check_10 = value_variable_222_to_check[11:6];
assign enable_variable_222_to_check_10 = enable_variable_222_to_check;

// 对校验节点107传递过来的数据进行整合
assign value_check_to_variable_222[17:12] = value_check_107_to_variable_222;
assign enable_check_to_variable_222[2] = enable_check_107_to_variable_222;
// 将变量节点222的输出与校验节点107的输入相连
assign value_variable_222_to_check_107 = value_variable_222_to_check[17:12];
assign enable_variable_222_to_check_107 = enable_variable_222_to_check;


// 变量节点223的接口
wire [17:0] value_check_to_variable_223;
wire [2:0] enable_check_to_variable_223;
wire [5:0] value_variable_223_to_decision;
wire [17:0] value_variable_223_to_check;

wire enable_variable_223_to_check;
// 对校验节点9传递过来的数据进行整合
assign value_check_to_variable_223[5:0] = value_check_9_to_variable_223;
assign enable_check_to_variable_223[0] = enable_check_9_to_variable_223;
// 将变量节点223的输出与校验节点9的输入相连
assign value_variable_223_to_check_9 = value_variable_223_to_check[5:0];
assign enable_variable_223_to_check_9 = enable_variable_223_to_check;

// 对校验节点67传递过来的数据进行整合
assign value_check_to_variable_223[11:6] = value_check_67_to_variable_223;
assign enable_check_to_variable_223[1] = enable_check_67_to_variable_223;
// 将变量节点223的输出与校验节点67的输入相连
assign value_variable_223_to_check_67 = value_variable_223_to_check[11:6];
assign enable_variable_223_to_check_67 = enable_variable_223_to_check;

// 对校验节点100传递过来的数据进行整合
assign value_check_to_variable_223[17:12] = value_check_100_to_variable_223;
assign enable_check_to_variable_223[2] = enable_check_100_to_variable_223;
// 将变量节点223的输出与校验节点100的输入相连
assign value_variable_223_to_check_100 = value_variable_223_to_check[17:12];
assign enable_variable_223_to_check_100 = enable_variable_223_to_check;


// 变量节点224的接口
wire [17:0] value_check_to_variable_224;
wire [2:0] enable_check_to_variable_224;
wire [5:0] value_variable_224_to_decision;
wire [17:0] value_variable_224_to_check;

wire enable_variable_224_to_check;
// 对校验节点11传递过来的数据进行整合
assign value_check_to_variable_224[5:0] = value_check_11_to_variable_224;
assign enable_check_to_variable_224[0] = enable_check_11_to_variable_224;
// 将变量节点224的输出与校验节点11的输入相连
assign value_variable_224_to_check_11 = value_variable_224_to_check[5:0];
assign enable_variable_224_to_check_11 = enable_variable_224_to_check;

// 对校验节点56传递过来的数据进行整合
assign value_check_to_variable_224[11:6] = value_check_56_to_variable_224;
assign enable_check_to_variable_224[1] = enable_check_56_to_variable_224;
// 将变量节点224的输出与校验节点56的输入相连
assign value_variable_224_to_check_56 = value_variable_224_to_check[11:6];
assign enable_variable_224_to_check_56 = enable_variable_224_to_check;

// 对校验节点116传递过来的数据进行整合
assign value_check_to_variable_224[17:12] = value_check_116_to_variable_224;
assign enable_check_to_variable_224[2] = enable_check_116_to_variable_224;
// 将变量节点224的输出与校验节点116的输入相连
assign value_variable_224_to_check_116 = value_variable_224_to_check[17:12];
assign enable_variable_224_to_check_116 = enable_variable_224_to_check;


// 变量节点225的接口
wire [17:0] value_check_to_variable_225;
wire [2:0] enable_check_to_variable_225;
wire [5:0] value_variable_225_to_decision;
wire [17:0] value_variable_225_to_check;

wire enable_variable_225_to_check;
// 对校验节点12传递过来的数据进行整合
assign value_check_to_variable_225[5:0] = value_check_12_to_variable_225;
assign enable_check_to_variable_225[0] = enable_check_12_to_variable_225;
// 将变量节点225的输出与校验节点12的输入相连
assign value_variable_225_to_check_12 = value_variable_225_to_check[5:0];
assign enable_variable_225_to_check_12 = enable_variable_225_to_check;

// 对校验节点27传递过来的数据进行整合
assign value_check_to_variable_225[11:6] = value_check_27_to_variable_225;
assign enable_check_to_variable_225[1] = enable_check_27_to_variable_225;
// 将变量节点225的输出与校验节点27的输入相连
assign value_variable_225_to_check_27 = value_variable_225_to_check[11:6];
assign enable_variable_225_to_check_27 = enable_variable_225_to_check;

// 对校验节点33传递过来的数据进行整合
assign value_check_to_variable_225[17:12] = value_check_33_to_variable_225;
assign enable_check_to_variable_225[2] = enable_check_33_to_variable_225;
// 将变量节点225的输出与校验节点33的输入相连
assign value_variable_225_to_check_33 = value_variable_225_to_check[17:12];
assign enable_variable_225_to_check_33 = enable_variable_225_to_check;


// 变量节点226的接口
wire [17:0] value_check_to_variable_226;
wire [2:0] enable_check_to_variable_226;
wire [5:0] value_variable_226_to_decision;
wire [17:0] value_variable_226_to_check;

wire enable_variable_226_to_check;
// 对校验节点13传递过来的数据进行整合
assign value_check_to_variable_226[5:0] = value_check_13_to_variable_226;
assign enable_check_to_variable_226[0] = enable_check_13_to_variable_226;
// 将变量节点226的输出与校验节点13的输入相连
assign value_variable_226_to_check_13 = value_variable_226_to_check[5:0];
assign enable_variable_226_to_check_13 = enable_variable_226_to_check;

// 对校验节点22传递过来的数据进行整合
assign value_check_to_variable_226[11:6] = value_check_22_to_variable_226;
assign enable_check_to_variable_226[1] = enable_check_22_to_variable_226;
// 将变量节点226的输出与校验节点22的输入相连
assign value_variable_226_to_check_22 = value_variable_226_to_check[11:6];
assign enable_variable_226_to_check_22 = enable_variable_226_to_check;

// 对校验节点92传递过来的数据进行整合
assign value_check_to_variable_226[17:12] = value_check_92_to_variable_226;
assign enable_check_to_variable_226[2] = enable_check_92_to_variable_226;
// 将变量节点226的输出与校验节点92的输入相连
assign value_variable_226_to_check_92 = value_variable_226_to_check[17:12];
assign enable_variable_226_to_check_92 = enable_variable_226_to_check;


// 变量节点227的接口
wire [17:0] value_check_to_variable_227;
wire [2:0] enable_check_to_variable_227;
wire [5:0] value_variable_227_to_decision;
wire [17:0] value_variable_227_to_check;

wire enable_variable_227_to_check;
// 对校验节点14传递过来的数据进行整合
assign value_check_to_variable_227[5:0] = value_check_14_to_variable_227;
assign enable_check_to_variable_227[0] = enable_check_14_to_variable_227;
// 将变量节点227的输出与校验节点14的输入相连
assign value_variable_227_to_check_14 = value_variable_227_to_check[5:0];
assign enable_variable_227_to_check_14 = enable_variable_227_to_check;

// 对校验节点45传递过来的数据进行整合
assign value_check_to_variable_227[11:6] = value_check_45_to_variable_227;
assign enable_check_to_variable_227[1] = enable_check_45_to_variable_227;
// 将变量节点227的输出与校验节点45的输入相连
assign value_variable_227_to_check_45 = value_variable_227_to_check[11:6];
assign enable_variable_227_to_check_45 = enable_variable_227_to_check;

// 对校验节点71传递过来的数据进行整合
assign value_check_to_variable_227[17:12] = value_check_71_to_variable_227;
assign enable_check_to_variable_227[2] = enable_check_71_to_variable_227;
// 将变量节点227的输出与校验节点71的输入相连
assign value_variable_227_to_check_71 = value_variable_227_to_check[17:12];
assign enable_variable_227_to_check_71 = enable_variable_227_to_check;


// 变量节点228的接口
wire [17:0] value_check_to_variable_228;
wire [2:0] enable_check_to_variable_228;
wire [5:0] value_variable_228_to_decision;
wire [17:0] value_variable_228_to_check;

wire enable_variable_228_to_check;
// 对校验节点17传递过来的数据进行整合
assign value_check_to_variable_228[5:0] = value_check_17_to_variable_228;
assign enable_check_to_variable_228[0] = enable_check_17_to_variable_228;
// 将变量节点228的输出与校验节点17的输入相连
assign value_variable_228_to_check_17 = value_variable_228_to_check[5:0];
assign enable_variable_228_to_check_17 = enable_variable_228_to_check;

// 对校验节点47传递过来的数据进行整合
assign value_check_to_variable_228[11:6] = value_check_47_to_variable_228;
assign enable_check_to_variable_228[1] = enable_check_47_to_variable_228;
// 将变量节点228的输出与校验节点47的输入相连
assign value_variable_228_to_check_47 = value_variable_228_to_check[11:6];
assign enable_variable_228_to_check_47 = enable_variable_228_to_check;

// 对校验节点57传递过来的数据进行整合
assign value_check_to_variable_228[17:12] = value_check_57_to_variable_228;
assign enable_check_to_variable_228[2] = enable_check_57_to_variable_228;
// 将变量节点228的输出与校验节点57的输入相连
assign value_variable_228_to_check_57 = value_variable_228_to_check[17:12];
assign enable_variable_228_to_check_57 = enable_variable_228_to_check;


// 变量节点229的接口
wire [17:0] value_check_to_variable_229;
wire [2:0] enable_check_to_variable_229;
wire [5:0] value_variable_229_to_decision;
wire [17:0] value_variable_229_to_check;

wire enable_variable_229_to_check;
// 对校验节点18传递过来的数据进行整合
assign value_check_to_variable_229[5:0] = value_check_18_to_variable_229;
assign enable_check_to_variable_229[0] = enable_check_18_to_variable_229;
// 将变量节点229的输出与校验节点18的输入相连
assign value_variable_229_to_check_18 = value_variable_229_to_check[5:0];
assign enable_variable_229_to_check_18 = enable_variable_229_to_check;

// 对校验节点34传递过来的数据进行整合
assign value_check_to_variable_229[11:6] = value_check_34_to_variable_229;
assign enable_check_to_variable_229[1] = enable_check_34_to_variable_229;
// 将变量节点229的输出与校验节点34的输入相连
assign value_variable_229_to_check_34 = value_variable_229_to_check[11:6];
assign enable_variable_229_to_check_34 = enable_variable_229_to_check;

// 对校验节点102传递过来的数据进行整合
assign value_check_to_variable_229[17:12] = value_check_102_to_variable_229;
assign enable_check_to_variable_229[2] = enable_check_102_to_variable_229;
// 将变量节点229的输出与校验节点102的输入相连
assign value_variable_229_to_check_102 = value_variable_229_to_check[17:12];
assign enable_variable_229_to_check_102 = enable_variable_229_to_check;


// 变量节点230的接口
wire [17:0] value_check_to_variable_230;
wire [2:0] enable_check_to_variable_230;
wire [5:0] value_variable_230_to_decision;
wire [17:0] value_variable_230_to_check;

wire enable_variable_230_to_check;
// 对校验节点19传递过来的数据进行整合
assign value_check_to_variable_230[5:0] = value_check_19_to_variable_230;
assign enable_check_to_variable_230[0] = enable_check_19_to_variable_230;
// 将变量节点230的输出与校验节点19的输入相连
assign value_variable_230_to_check_19 = value_variable_230_to_check[5:0];
assign enable_variable_230_to_check_19 = enable_variable_230_to_check;

// 对校验节点35传递过来的数据进行整合
assign value_check_to_variable_230[11:6] = value_check_35_to_variable_230;
assign enable_check_to_variable_230[1] = enable_check_35_to_variable_230;
// 将变量节点230的输出与校验节点35的输入相连
assign value_variable_230_to_check_35 = value_variable_230_to_check[11:6];
assign enable_variable_230_to_check_35 = enable_variable_230_to_check;

// 对校验节点91传递过来的数据进行整合
assign value_check_to_variable_230[17:12] = value_check_91_to_variable_230;
assign enable_check_to_variable_230[2] = enable_check_91_to_variable_230;
// 将变量节点230的输出与校验节点91的输入相连
assign value_variable_230_to_check_91 = value_variable_230_to_check[17:12];
assign enable_variable_230_to_check_91 = enable_variable_230_to_check;


// 变量节点231的接口
wire [17:0] value_check_to_variable_231;
wire [2:0] enable_check_to_variable_231;
wire [5:0] value_variable_231_to_decision;
wire [17:0] value_variable_231_to_check;

wire enable_variable_231_to_check;
// 对校验节点20传递过来的数据进行整合
assign value_check_to_variable_231[5:0] = value_check_20_to_variable_231;
assign enable_check_to_variable_231[0] = enable_check_20_to_variable_231;
// 将变量节点231的输出与校验节点20的输入相连
assign value_variable_231_to_check_20 = value_variable_231_to_check[5:0];
assign enable_variable_231_to_check_20 = enable_variable_231_to_check;

// 对校验节点44传递过来的数据进行整合
assign value_check_to_variable_231[11:6] = value_check_44_to_variable_231;
assign enable_check_to_variable_231[1] = enable_check_44_to_variable_231;
// 将变量节点231的输出与校验节点44的输入相连
assign value_variable_231_to_check_44 = value_variable_231_to_check[11:6];
assign enable_variable_231_to_check_44 = enable_variable_231_to_check;

// 对校验节点52传递过来的数据进行整合
assign value_check_to_variable_231[17:12] = value_check_52_to_variable_231;
assign enable_check_to_variable_231[2] = enable_check_52_to_variable_231;
// 将变量节点231的输出与校验节点52的输入相连
assign value_variable_231_to_check_52 = value_variable_231_to_check[17:12];
assign enable_variable_231_to_check_52 = enable_variable_231_to_check;


// 变量节点232的接口
wire [17:0] value_check_to_variable_232;
wire [2:0] enable_check_to_variable_232;
wire [5:0] value_variable_232_to_decision;
wire [17:0] value_variable_232_to_check;

wire enable_variable_232_to_check;
// 对校验节点23传递过来的数据进行整合
assign value_check_to_variable_232[5:0] = value_check_23_to_variable_232;
assign enable_check_to_variable_232[0] = enable_check_23_to_variable_232;
// 将变量节点232的输出与校验节点23的输入相连
assign value_variable_232_to_check_23 = value_variable_232_to_check[5:0];
assign enable_variable_232_to_check_23 = enable_variable_232_to_check;

// 对校验节点42传递过来的数据进行整合
assign value_check_to_variable_232[11:6] = value_check_42_to_variable_232;
assign enable_check_to_variable_232[1] = enable_check_42_to_variable_232;
// 将变量节点232的输出与校验节点42的输入相连
assign value_variable_232_to_check_42 = value_variable_232_to_check[11:6];
assign enable_variable_232_to_check_42 = enable_variable_232_to_check;

// 对校验节点86传递过来的数据进行整合
assign value_check_to_variable_232[17:12] = value_check_86_to_variable_232;
assign enable_check_to_variable_232[2] = enable_check_86_to_variable_232;
// 将变量节点232的输出与校验节点86的输入相连
assign value_variable_232_to_check_86 = value_variable_232_to_check[17:12];
assign enable_variable_232_to_check_86 = enable_variable_232_to_check;


// 变量节点233的接口
wire [17:0] value_check_to_variable_233;
wire [2:0] enable_check_to_variable_233;
wire [5:0] value_variable_233_to_decision;
wire [17:0] value_variable_233_to_check;

wire enable_variable_233_to_check;
// 对校验节点24传递过来的数据进行整合
assign value_check_to_variable_233[5:0] = value_check_24_to_variable_233;
assign enable_check_to_variable_233[0] = enable_check_24_to_variable_233;
// 将变量节点233的输出与校验节点24的输入相连
assign value_variable_233_to_check_24 = value_variable_233_to_check[5:0];
assign enable_variable_233_to_check_24 = enable_variable_233_to_check;

// 对校验节点54传递过来的数据进行整合
assign value_check_to_variable_233[11:6] = value_check_54_to_variable_233;
assign enable_check_to_variable_233[1] = enable_check_54_to_variable_233;
// 将变量节点233的输出与校验节点54的输入相连
assign value_variable_233_to_check_54 = value_variable_233_to_check[11:6];
assign enable_variable_233_to_check_54 = enable_variable_233_to_check;

// 对校验节点98传递过来的数据进行整合
assign value_check_to_variable_233[17:12] = value_check_98_to_variable_233;
assign enable_check_to_variable_233[2] = enable_check_98_to_variable_233;
// 将变量节点233的输出与校验节点98的输入相连
assign value_variable_233_to_check_98 = value_variable_233_to_check[17:12];
assign enable_variable_233_to_check_98 = enable_variable_233_to_check;


// 变量节点234的接口
wire [17:0] value_check_to_variable_234;
wire [2:0] enable_check_to_variable_234;
wire [5:0] value_variable_234_to_decision;
wire [17:0] value_variable_234_to_check;

wire enable_variable_234_to_check;
// 对校验节点25传递过来的数据进行整合
assign value_check_to_variable_234[5:0] = value_check_25_to_variable_234;
assign enable_check_to_variable_234[0] = enable_check_25_to_variable_234;
// 将变量节点234的输出与校验节点25的输入相连
assign value_variable_234_to_check_25 = value_variable_234_to_check[5:0];
assign enable_variable_234_to_check_25 = enable_variable_234_to_check;

// 对校验节点75传递过来的数据进行整合
assign value_check_to_variable_234[11:6] = value_check_75_to_variable_234;
assign enable_check_to_variable_234[1] = enable_check_75_to_variable_234;
// 将变量节点234的输出与校验节点75的输入相连
assign value_variable_234_to_check_75 = value_variable_234_to_check[11:6];
assign enable_variable_234_to_check_75 = enable_variable_234_to_check;

// 对校验节点81传递过来的数据进行整合
assign value_check_to_variable_234[17:12] = value_check_81_to_variable_234;
assign enable_check_to_variable_234[2] = enable_check_81_to_variable_234;
// 将变量节点234的输出与校验节点81的输入相连
assign value_variable_234_to_check_81 = value_variable_234_to_check[17:12];
assign enable_variable_234_to_check_81 = enable_variable_234_to_check;


// 变量节点235的接口
wire [17:0] value_check_to_variable_235;
wire [2:0] enable_check_to_variable_235;
wire [5:0] value_variable_235_to_decision;
wire [17:0] value_variable_235_to_check;

wire enable_variable_235_to_check;
// 对校验节点26传递过来的数据进行整合
assign value_check_to_variable_235[5:0] = value_check_26_to_variable_235;
assign enable_check_to_variable_235[0] = enable_check_26_to_variable_235;
// 将变量节点235的输出与校验节点26的输入相连
assign value_variable_235_to_check_26 = value_variable_235_to_check[5:0];
assign enable_variable_235_to_check_26 = enable_variable_235_to_check;

// 对校验节点50传递过来的数据进行整合
assign value_check_to_variable_235[11:6] = value_check_50_to_variable_235;
assign enable_check_to_variable_235[1] = enable_check_50_to_variable_235;
// 将变量节点235的输出与校验节点50的输入相连
assign value_variable_235_to_check_50 = value_variable_235_to_check[11:6];
assign enable_variable_235_to_check_50 = enable_variable_235_to_check;

// 对校验节点125传递过来的数据进行整合
assign value_check_to_variable_235[17:12] = value_check_125_to_variable_235;
assign enable_check_to_variable_235[2] = enable_check_125_to_variable_235;
// 将变量节点235的输出与校验节点125的输入相连
assign value_variable_235_to_check_125 = value_variable_235_to_check[17:12];
assign enable_variable_235_to_check_125 = enable_variable_235_to_check;


// 变量节点236的接口
wire [17:0] value_check_to_variable_236;
wire [2:0] enable_check_to_variable_236;
wire [5:0] value_variable_236_to_decision;
wire [17:0] value_variable_236_to_check;

wire enable_variable_236_to_check;
// 对校验节点28传递过来的数据进行整合
assign value_check_to_variable_236[5:0] = value_check_28_to_variable_236;
assign enable_check_to_variable_236[0] = enable_check_28_to_variable_236;
// 将变量节点236的输出与校验节点28的输入相连
assign value_variable_236_to_check_28 = value_variable_236_to_check[5:0];
assign enable_variable_236_to_check_28 = enable_variable_236_to_check;

// 对校验节点31传递过来的数据进行整合
assign value_check_to_variable_236[11:6] = value_check_31_to_variable_236;
assign enable_check_to_variable_236[1] = enable_check_31_to_variable_236;
// 将变量节点236的输出与校验节点31的输入相连
assign value_variable_236_to_check_31 = value_variable_236_to_check[11:6];
assign enable_variable_236_to_check_31 = enable_variable_236_to_check;

// 对校验节点109传递过来的数据进行整合
assign value_check_to_variable_236[17:12] = value_check_109_to_variable_236;
assign enable_check_to_variable_236[2] = enable_check_109_to_variable_236;
// 将变量节点236的输出与校验节点109的输入相连
assign value_variable_236_to_check_109 = value_variable_236_to_check[17:12];
assign enable_variable_236_to_check_109 = enable_variable_236_to_check;


// 变量节点237的接口
wire [17:0] value_check_to_variable_237;
wire [2:0] enable_check_to_variable_237;
wire [5:0] value_variable_237_to_decision;
wire [17:0] value_variable_237_to_check;

wire enable_variable_237_to_check;
// 对校验节点29传递过来的数据进行整合
assign value_check_to_variable_237[5:0] = value_check_29_to_variable_237;
assign enable_check_to_variable_237[0] = enable_check_29_to_variable_237;
// 将变量节点237的输出与校验节点29的输入相连
assign value_variable_237_to_check_29 = value_variable_237_to_check[5:0];
assign enable_variable_237_to_check_29 = enable_variable_237_to_check;

// 对校验节点104传递过来的数据进行整合
assign value_check_to_variable_237[11:6] = value_check_104_to_variable_237;
assign enable_check_to_variable_237[1] = enable_check_104_to_variable_237;
// 将变量节点237的输出与校验节点104的输入相连
assign value_variable_237_to_check_104 = value_variable_237_to_check[11:6];
assign enable_variable_237_to_check_104 = enable_variable_237_to_check;

// 对校验节点121传递过来的数据进行整合
assign value_check_to_variable_237[17:12] = value_check_121_to_variable_237;
assign enable_check_to_variable_237[2] = enable_check_121_to_variable_237;
// 将变量节点237的输出与校验节点121的输入相连
assign value_variable_237_to_check_121 = value_variable_237_to_check[17:12];
assign enable_variable_237_to_check_121 = enable_variable_237_to_check;


// 变量节点238的接口
wire [17:0] value_check_to_variable_238;
wire [2:0] enable_check_to_variable_238;
wire [5:0] value_variable_238_to_decision;
wire [17:0] value_variable_238_to_check;

wire enable_variable_238_to_check;
// 对校验节点36传递过来的数据进行整合
assign value_check_to_variable_238[5:0] = value_check_36_to_variable_238;
assign enable_check_to_variable_238[0] = enable_check_36_to_variable_238;
// 将变量节点238的输出与校验节点36的输入相连
assign value_variable_238_to_check_36 = value_variable_238_to_check[5:0];
assign enable_variable_238_to_check_36 = enable_variable_238_to_check;

// 对校验节点113传递过来的数据进行整合
assign value_check_to_variable_238[11:6] = value_check_113_to_variable_238;
assign enable_check_to_variable_238[1] = enable_check_113_to_variable_238;
// 将变量节点238的输出与校验节点113的输入相连
assign value_variable_238_to_check_113 = value_variable_238_to_check[11:6];
assign enable_variable_238_to_check_113 = enable_variable_238_to_check;

// 对校验节点120传递过来的数据进行整合
assign value_check_to_variable_238[17:12] = value_check_120_to_variable_238;
assign enable_check_to_variable_238[2] = enable_check_120_to_variable_238;
// 将变量节点238的输出与校验节点120的输入相连
assign value_variable_238_to_check_120 = value_variable_238_to_check[17:12];
assign enable_variable_238_to_check_120 = enable_variable_238_to_check;


// 变量节点239的接口
wire [17:0] value_check_to_variable_239;
wire [2:0] enable_check_to_variable_239;
wire [5:0] value_variable_239_to_decision;
wire [17:0] value_variable_239_to_check;

wire enable_variable_239_to_check;
// 对校验节点39传递过来的数据进行整合
assign value_check_to_variable_239[5:0] = value_check_39_to_variable_239;
assign enable_check_to_variable_239[0] = enable_check_39_to_variable_239;
// 将变量节点239的输出与校验节点39的输入相连
assign value_variable_239_to_check_39 = value_variable_239_to_check[5:0];
assign enable_variable_239_to_check_39 = enable_variable_239_to_check;

// 对校验节点64传递过来的数据进行整合
assign value_check_to_variable_239[11:6] = value_check_64_to_variable_239;
assign enable_check_to_variable_239[1] = enable_check_64_to_variable_239;
// 将变量节点239的输出与校验节点64的输入相连
assign value_variable_239_to_check_64 = value_variable_239_to_check[11:6];
assign enable_variable_239_to_check_64 = enable_variable_239_to_check;

// 对校验节点87传递过来的数据进行整合
assign value_check_to_variable_239[17:12] = value_check_87_to_variable_239;
assign enable_check_to_variable_239[2] = enable_check_87_to_variable_239;
// 将变量节点239的输出与校验节点87的输入相连
assign value_variable_239_to_check_87 = value_variable_239_to_check[17:12];
assign enable_variable_239_to_check_87 = enable_variable_239_to_check;


// 变量节点240的接口
wire [17:0] value_check_to_variable_240;
wire [2:0] enable_check_to_variable_240;
wire [5:0] value_variable_240_to_decision;
wire [17:0] value_variable_240_to_check;

wire enable_variable_240_to_check;
// 对校验节点40传递过来的数据进行整合
assign value_check_to_variable_240[5:0] = value_check_40_to_variable_240;
assign enable_check_to_variable_240[0] = enable_check_40_to_variable_240;
// 将变量节点240的输出与校验节点40的输入相连
assign value_variable_240_to_check_40 = value_variable_240_to_check[5:0];
assign enable_variable_240_to_check_40 = enable_variable_240_to_check;

// 对校验节点49传递过来的数据进行整合
assign value_check_to_variable_240[11:6] = value_check_49_to_variable_240;
assign enable_check_to_variable_240[1] = enable_check_49_to_variable_240;
// 将变量节点240的输出与校验节点49的输入相连
assign value_variable_240_to_check_49 = value_variable_240_to_check[11:6];
assign enable_variable_240_to_check_49 = enable_variable_240_to_check;

// 对校验节点97传递过来的数据进行整合
assign value_check_to_variable_240[17:12] = value_check_97_to_variable_240;
assign enable_check_to_variable_240[2] = enable_check_97_to_variable_240;
// 将变量节点240的输出与校验节点97的输入相连
assign value_variable_240_to_check_97 = value_variable_240_to_check[17:12];
assign enable_variable_240_to_check_97 = enable_variable_240_to_check;


// 变量节点241的接口
wire [17:0] value_check_to_variable_241;
wire [2:0] enable_check_to_variable_241;
wire [5:0] value_variable_241_to_decision;
wire [17:0] value_variable_241_to_check;

wire enable_variable_241_to_check;
// 对校验节点41传递过来的数据进行整合
assign value_check_to_variable_241[5:0] = value_check_41_to_variable_241;
assign enable_check_to_variable_241[0] = enable_check_41_to_variable_241;
// 将变量节点241的输出与校验节点41的输入相连
assign value_variable_241_to_check_41 = value_variable_241_to_check[5:0];
assign enable_variable_241_to_check_41 = enable_variable_241_to_check;

// 对校验节点110传递过来的数据进行整合
assign value_check_to_variable_241[11:6] = value_check_110_to_variable_241;
assign enable_check_to_variable_241[1] = enable_check_110_to_variable_241;
// 将变量节点241的输出与校验节点110的输入相连
assign value_variable_241_to_check_110 = value_variable_241_to_check[11:6];
assign enable_variable_241_to_check_110 = enable_variable_241_to_check;

// 对校验节点112传递过来的数据进行整合
assign value_check_to_variable_241[17:12] = value_check_112_to_variable_241;
assign enable_check_to_variable_241[2] = enable_check_112_to_variable_241;
// 将变量节点241的输出与校验节点112的输入相连
assign value_variable_241_to_check_112 = value_variable_241_to_check[17:12];
assign enable_variable_241_to_check_112 = enable_variable_241_to_check;


// 变量节点242的接口
wire [17:0] value_check_to_variable_242;
wire [2:0] enable_check_to_variable_242;
wire [5:0] value_variable_242_to_decision;
wire [17:0] value_variable_242_to_check;

wire enable_variable_242_to_check;
// 对校验节点46传递过来的数据进行整合
assign value_check_to_variable_242[5:0] = value_check_46_to_variable_242;
assign enable_check_to_variable_242[0] = enable_check_46_to_variable_242;
// 将变量节点242的输出与校验节点46的输入相连
assign value_variable_242_to_check_46 = value_variable_242_to_check[5:0];
assign enable_variable_242_to_check_46 = enable_variable_242_to_check;

// 对校验节点61传递过来的数据进行整合
assign value_check_to_variable_242[11:6] = value_check_61_to_variable_242;
assign enable_check_to_variable_242[1] = enable_check_61_to_variable_242;
// 将变量节点242的输出与校验节点61的输入相连
assign value_variable_242_to_check_61 = value_variable_242_to_check[11:6];
assign enable_variable_242_to_check_61 = enable_variable_242_to_check;

// 对校验节点79传递过来的数据进行整合
assign value_check_to_variable_242[17:12] = value_check_79_to_variable_242;
assign enable_check_to_variable_242[2] = enable_check_79_to_variable_242;
// 将变量节点242的输出与校验节点79的输入相连
assign value_variable_242_to_check_79 = value_variable_242_to_check[17:12];
assign enable_variable_242_to_check_79 = enable_variable_242_to_check;


// 变量节点243的接口
wire [17:0] value_check_to_variable_243;
wire [2:0] enable_check_to_variable_243;
wire [5:0] value_variable_243_to_decision;
wire [17:0] value_variable_243_to_check;

wire enable_variable_243_to_check;
// 对校验节点48传递过来的数据进行整合
assign value_check_to_variable_243[5:0] = value_check_48_to_variable_243;
assign enable_check_to_variable_243[0] = enable_check_48_to_variable_243;
// 将变量节点243的输出与校验节点48的输入相连
assign value_variable_243_to_check_48 = value_variable_243_to_check[5:0];
assign enable_variable_243_to_check_48 = enable_variable_243_to_check;

// 对校验节点53传递过来的数据进行整合
assign value_check_to_variable_243[11:6] = value_check_53_to_variable_243;
assign enable_check_to_variable_243[1] = enable_check_53_to_variable_243;
// 将变量节点243的输出与校验节点53的输入相连
assign value_variable_243_to_check_53 = value_variable_243_to_check[11:6];
assign enable_variable_243_to_check_53 = enable_variable_243_to_check;

// 对校验节点84传递过来的数据进行整合
assign value_check_to_variable_243[17:12] = value_check_84_to_variable_243;
assign enable_check_to_variable_243[2] = enable_check_84_to_variable_243;
// 将变量节点243的输出与校验节点84的输入相连
assign value_variable_243_to_check_84 = value_variable_243_to_check[17:12];
assign enable_variable_243_to_check_84 = enable_variable_243_to_check;


// 变量节点244的接口
wire [17:0] value_check_to_variable_244;
wire [2:0] enable_check_to_variable_244;
wire [5:0] value_variable_244_to_decision;
wire [17:0] value_variable_244_to_check;

wire enable_variable_244_to_check;
// 对校验节点51传递过来的数据进行整合
assign value_check_to_variable_244[5:0] = value_check_51_to_variable_244;
assign enable_check_to_variable_244[0] = enable_check_51_to_variable_244;
// 将变量节点244的输出与校验节点51的输入相连
assign value_variable_244_to_check_51 = value_variable_244_to_check[5:0];
assign enable_variable_244_to_check_51 = enable_variable_244_to_check;

// 对校验节点94传递过来的数据进行整合
assign value_check_to_variable_244[11:6] = value_check_94_to_variable_244;
assign enable_check_to_variable_244[1] = enable_check_94_to_variable_244;
// 将变量节点244的输出与校验节点94的输入相连
assign value_variable_244_to_check_94 = value_variable_244_to_check[11:6];
assign enable_variable_244_to_check_94 = enable_variable_244_to_check;

// 对校验节点126传递过来的数据进行整合
assign value_check_to_variable_244[17:12] = value_check_126_to_variable_244;
assign enable_check_to_variable_244[2] = enable_check_126_to_variable_244;
// 将变量节点244的输出与校验节点126的输入相连
assign value_variable_244_to_check_126 = value_variable_244_to_check[17:12];
assign enable_variable_244_to_check_126 = enable_variable_244_to_check;


// 变量节点245的接口
wire [17:0] value_check_to_variable_245;
wire [2:0] enable_check_to_variable_245;
wire [5:0] value_variable_245_to_decision;
wire [17:0] value_variable_245_to_check;

wire enable_variable_245_to_check;
// 对校验节点55传递过来的数据进行整合
assign value_check_to_variable_245[5:0] = value_check_55_to_variable_245;
assign enable_check_to_variable_245[0] = enable_check_55_to_variable_245;
// 将变量节点245的输出与校验节点55的输入相连
assign value_variable_245_to_check_55 = value_variable_245_to_check[5:0];
assign enable_variable_245_to_check_55 = enable_variable_245_to_check;

// 对校验节点77传递过来的数据进行整合
assign value_check_to_variable_245[11:6] = value_check_77_to_variable_245;
assign enable_check_to_variable_245[1] = enable_check_77_to_variable_245;
// 将变量节点245的输出与校验节点77的输入相连
assign value_variable_245_to_check_77 = value_variable_245_to_check[11:6];
assign enable_variable_245_to_check_77 = enable_variable_245_to_check;

// 对校验节点123传递过来的数据进行整合
assign value_check_to_variable_245[17:12] = value_check_123_to_variable_245;
assign enable_check_to_variable_245[2] = enable_check_123_to_variable_245;
// 将变量节点245的输出与校验节点123的输入相连
assign value_variable_245_to_check_123 = value_variable_245_to_check[17:12];
assign enable_variable_245_to_check_123 = enable_variable_245_to_check;


// 变量节点246的接口
wire [17:0] value_check_to_variable_246;
wire [2:0] enable_check_to_variable_246;
wire [5:0] value_variable_246_to_decision;
wire [17:0] value_variable_246_to_check;

wire enable_variable_246_to_check;
// 对校验节点58传递过来的数据进行整合
assign value_check_to_variable_246[5:0] = value_check_58_to_variable_246;
assign enable_check_to_variable_246[0] = enable_check_58_to_variable_246;
// 将变量节点246的输出与校验节点58的输入相连
assign value_variable_246_to_check_58 = value_variable_246_to_check[5:0];
assign enable_variable_246_to_check_58 = enable_variable_246_to_check;

// 对校验节点59传递过来的数据进行整合
assign value_check_to_variable_246[11:6] = value_check_59_to_variable_246;
assign enable_check_to_variable_246[1] = enable_check_59_to_variable_246;
// 将变量节点246的输出与校验节点59的输入相连
assign value_variable_246_to_check_59 = value_variable_246_to_check[11:6];
assign enable_variable_246_to_check_59 = enable_variable_246_to_check;

// 对校验节点90传递过来的数据进行整合
assign value_check_to_variable_246[17:12] = value_check_90_to_variable_246;
assign enable_check_to_variable_246[2] = enable_check_90_to_variable_246;
// 将变量节点246的输出与校验节点90的输入相连
assign value_variable_246_to_check_90 = value_variable_246_to_check[17:12];
assign enable_variable_246_to_check_90 = enable_variable_246_to_check;


// 变量节点247的接口
wire [17:0] value_check_to_variable_247;
wire [2:0] enable_check_to_variable_247;
wire [5:0] value_variable_247_to_decision;
wire [17:0] value_variable_247_to_check;

wire enable_variable_247_to_check;
// 对校验节点60传递过来的数据进行整合
assign value_check_to_variable_247[5:0] = value_check_60_to_variable_247;
assign enable_check_to_variable_247[0] = enable_check_60_to_variable_247;
// 将变量节点247的输出与校验节点60的输入相连
assign value_variable_247_to_check_60 = value_variable_247_to_check[5:0];
assign enable_variable_247_to_check_60 = enable_variable_247_to_check;

// 对校验节点88传递过来的数据进行整合
assign value_check_to_variable_247[11:6] = value_check_88_to_variable_247;
assign enable_check_to_variable_247[1] = enable_check_88_to_variable_247;
// 将变量节点247的输出与校验节点88的输入相连
assign value_variable_247_to_check_88 = value_variable_247_to_check[11:6];
assign enable_variable_247_to_check_88 = enable_variable_247_to_check;

// 对校验节点93传递过来的数据进行整合
assign value_check_to_variable_247[17:12] = value_check_93_to_variable_247;
assign enable_check_to_variable_247[2] = enable_check_93_to_variable_247;
// 将变量节点247的输出与校验节点93的输入相连
assign value_variable_247_to_check_93 = value_variable_247_to_check[17:12];
assign enable_variable_247_to_check_93 = enable_variable_247_to_check;


// 变量节点248的接口
wire [17:0] value_check_to_variable_248;
wire [2:0] enable_check_to_variable_248;
wire [5:0] value_variable_248_to_decision;
wire [17:0] value_variable_248_to_check;

wire enable_variable_248_to_check;
// 对校验节点62传递过来的数据进行整合
assign value_check_to_variable_248[5:0] = value_check_62_to_variable_248;
assign enable_check_to_variable_248[0] = enable_check_62_to_variable_248;
// 将变量节点248的输出与校验节点62的输入相连
assign value_variable_248_to_check_62 = value_variable_248_to_check[5:0];
assign enable_variable_248_to_check_62 = enable_variable_248_to_check;

// 对校验节点66传递过来的数据进行整合
assign value_check_to_variable_248[11:6] = value_check_66_to_variable_248;
assign enable_check_to_variable_248[1] = enable_check_66_to_variable_248;
// 将变量节点248的输出与校验节点66的输入相连
assign value_variable_248_to_check_66 = value_variable_248_to_check[11:6];
assign enable_variable_248_to_check_66 = enable_variable_248_to_check;

// 对校验节点124传递过来的数据进行整合
assign value_check_to_variable_248[17:12] = value_check_124_to_variable_248;
assign enable_check_to_variable_248[2] = enable_check_124_to_variable_248;
// 将变量节点248的输出与校验节点124的输入相连
assign value_variable_248_to_check_124 = value_variable_248_to_check[17:12];
assign enable_variable_248_to_check_124 = enable_variable_248_to_check;


// 变量节点249的接口
wire [17:0] value_check_to_variable_249;
wire [2:0] enable_check_to_variable_249;
wire [5:0] value_variable_249_to_decision;
wire [17:0] value_variable_249_to_check;

wire enable_variable_249_to_check;
// 对校验节点65传递过来的数据进行整合
assign value_check_to_variable_249[5:0] = value_check_65_to_variable_249;
assign enable_check_to_variable_249[0] = enable_check_65_to_variable_249;
// 将变量节点249的输出与校验节点65的输入相连
assign value_variable_249_to_check_65 = value_variable_249_to_check[5:0];
assign enable_variable_249_to_check_65 = enable_variable_249_to_check;

// 对校验节点74传递过来的数据进行整合
assign value_check_to_variable_249[11:6] = value_check_74_to_variable_249;
assign enable_check_to_variable_249[1] = enable_check_74_to_variable_249;
// 将变量节点249的输出与校验节点74的输入相连
assign value_variable_249_to_check_74 = value_variable_249_to_check[11:6];
assign enable_variable_249_to_check_74 = enable_variable_249_to_check;

// 对校验节点105传递过来的数据进行整合
assign value_check_to_variable_249[17:12] = value_check_105_to_variable_249;
assign enable_check_to_variable_249[2] = enable_check_105_to_variable_249;
// 将变量节点249的输出与校验节点105的输入相连
assign value_variable_249_to_check_105 = value_variable_249_to_check[17:12];
assign enable_variable_249_to_check_105 = enable_variable_249_to_check;


// 变量节点250的接口
wire [17:0] value_check_to_variable_250;
wire [2:0] enable_check_to_variable_250;
wire [5:0] value_variable_250_to_decision;
wire [17:0] value_variable_250_to_check;

wire enable_variable_250_to_check;
// 对校验节点68传递过来的数据进行整合
assign value_check_to_variable_250[5:0] = value_check_68_to_variable_250;
assign enable_check_to_variable_250[0] = enable_check_68_to_variable_250;
// 将变量节点250的输出与校验节点68的输入相连
assign value_variable_250_to_check_68 = value_variable_250_to_check[5:0];
assign enable_variable_250_to_check_68 = enable_variable_250_to_check;

// 对校验节点85传递过来的数据进行整合
assign value_check_to_variable_250[11:6] = value_check_85_to_variable_250;
assign enable_check_to_variable_250[1] = enable_check_85_to_variable_250;
// 将变量节点250的输出与校验节点85的输入相连
assign value_variable_250_to_check_85 = value_variable_250_to_check[11:6];
assign enable_variable_250_to_check_85 = enable_variable_250_to_check;

// 对校验节点96传递过来的数据进行整合
assign value_check_to_variable_250[17:12] = value_check_96_to_variable_250;
assign enable_check_to_variable_250[2] = enable_check_96_to_variable_250;
// 将变量节点250的输出与校验节点96的输入相连
assign value_variable_250_to_check_96 = value_variable_250_to_check[17:12];
assign enable_variable_250_to_check_96 = enable_variable_250_to_check;


// 变量节点251的接口
wire [17:0] value_check_to_variable_251;
wire [2:0] enable_check_to_variable_251;
wire [5:0] value_variable_251_to_decision;
wire [17:0] value_variable_251_to_check;

wire enable_variable_251_to_check;
// 对校验节点70传递过来的数据进行整合
assign value_check_to_variable_251[5:0] = value_check_70_to_variable_251;
assign enable_check_to_variable_251[0] = enable_check_70_to_variable_251;
// 将变量节点251的输出与校验节点70的输入相连
assign value_variable_251_to_check_70 = value_variable_251_to_check[5:0];
assign enable_variable_251_to_check_70 = enable_variable_251_to_check;

// 对校验节点103传递过来的数据进行整合
assign value_check_to_variable_251[11:6] = value_check_103_to_variable_251;
assign enable_check_to_variable_251[1] = enable_check_103_to_variable_251;
// 将变量节点251的输出与校验节点103的输入相连
assign value_variable_251_to_check_103 = value_variable_251_to_check[11:6];
assign enable_variable_251_to_check_103 = enable_variable_251_to_check;

// 对校验节点115传递过来的数据进行整合
assign value_check_to_variable_251[17:12] = value_check_115_to_variable_251;
assign enable_check_to_variable_251[2] = enable_check_115_to_variable_251;
// 将变量节点251的输出与校验节点115的输入相连
assign value_variable_251_to_check_115 = value_variable_251_to_check[17:12];
assign enable_variable_251_to_check_115 = enable_variable_251_to_check;


// 变量节点252的接口
wire [17:0] value_check_to_variable_252;
wire [2:0] enable_check_to_variable_252;
wire [5:0] value_variable_252_to_decision;
wire [17:0] value_variable_252_to_check;

wire enable_variable_252_to_check;
// 对校验节点72传递过来的数据进行整合
assign value_check_to_variable_252[5:0] = value_check_72_to_variable_252;
assign enable_check_to_variable_252[0] = enable_check_72_to_variable_252;
// 将变量节点252的输出与校验节点72的输入相连
assign value_variable_252_to_check_72 = value_variable_252_to_check[5:0];
assign enable_variable_252_to_check_72 = enable_variable_252_to_check;

// 对校验节点82传递过来的数据进行整合
assign value_check_to_variable_252[11:6] = value_check_82_to_variable_252;
assign enable_check_to_variable_252[1] = enable_check_82_to_variable_252;
// 将变量节点252的输出与校验节点82的输入相连
assign value_variable_252_to_check_82 = value_variable_252_to_check[11:6];
assign enable_variable_252_to_check_82 = enable_variable_252_to_check;

// 对校验节点118传递过来的数据进行整合
assign value_check_to_variable_252[17:12] = value_check_118_to_variable_252;
assign enable_check_to_variable_252[2] = enable_check_118_to_variable_252;
// 将变量节点252的输出与校验节点118的输入相连
assign value_variable_252_to_check_118 = value_variable_252_to_check[17:12];
assign enable_variable_252_to_check_118 = enable_variable_252_to_check;


// 变量节点253的接口
wire [17:0] value_check_to_variable_253;
wire [2:0] enable_check_to_variable_253;
wire [5:0] value_variable_253_to_decision;
wire [17:0] value_variable_253_to_check;

wire enable_variable_253_to_check;
// 对校验节点76传递过来的数据进行整合
assign value_check_to_variable_253[5:0] = value_check_76_to_variable_253;
assign enable_check_to_variable_253[0] = enable_check_76_to_variable_253;
// 将变量节点253的输出与校验节点76的输入相连
assign value_variable_253_to_check_76 = value_variable_253_to_check[5:0];
assign enable_variable_253_to_check_76 = enable_variable_253_to_check;

// 对校验节点108传递过来的数据进行整合
assign value_check_to_variable_253[11:6] = value_check_108_to_variable_253;
assign enable_check_to_variable_253[1] = enable_check_108_to_variable_253;
// 将变量节点253的输出与校验节点108的输入相连
assign value_variable_253_to_check_108 = value_variable_253_to_check[11:6];
assign enable_variable_253_to_check_108 = enable_variable_253_to_check;

// 对校验节点114传递过来的数据进行整合
assign value_check_to_variable_253[17:12] = value_check_114_to_variable_253;
assign enable_check_to_variable_253[2] = enable_check_114_to_variable_253;
// 将变量节点253的输出与校验节点114的输入相连
assign value_variable_253_to_check_114 = value_variable_253_to_check[17:12];
assign enable_variable_253_to_check_114 = enable_variable_253_to_check;


// 变量节点254的接口
wire [17:0] value_check_to_variable_254;
wire [2:0] enable_check_to_variable_254;
wire [5:0] value_variable_254_to_decision;
wire [17:0] value_variable_254_to_check;

wire enable_variable_254_to_check;
// 对校验节点80传递过来的数据进行整合
assign value_check_to_variable_254[5:0] = value_check_80_to_variable_254;
assign enable_check_to_variable_254[0] = enable_check_80_to_variable_254;
// 将变量节点254的输出与校验节点80的输入相连
assign value_variable_254_to_check_80 = value_variable_254_to_check[5:0];
assign enable_variable_254_to_check_80 = enable_variable_254_to_check;

// 对校验节点106传递过来的数据进行整合
assign value_check_to_variable_254[11:6] = value_check_106_to_variable_254;
assign enable_check_to_variable_254[1] = enable_check_106_to_variable_254;
// 将变量节点254的输出与校验节点106的输入相连
assign value_variable_254_to_check_106 = value_variable_254_to_check[11:6];
assign enable_variable_254_to_check_106 = enable_variable_254_to_check;

// 对校验节点127传递过来的数据进行整合
assign value_check_to_variable_254[17:12] = value_check_127_to_variable_254;
assign enable_check_to_variable_254[2] = enable_check_127_to_variable_254;
// 将变量节点254的输出与校验节点127的输入相连
assign value_variable_254_to_check_127 = value_variable_254_to_check[17:12];
assign enable_variable_254_to_check_127 = enable_variable_254_to_check;


// 变量节点255的接口
wire [17:0] value_check_to_variable_255;
wire [2:0] enable_check_to_variable_255;
wire [5:0] value_variable_255_to_decision;
wire [17:0] value_variable_255_to_check;

wire enable_variable_255_to_check;
// 对校验节点95传递过来的数据进行整合
assign value_check_to_variable_255[5:0] = value_check_95_to_variable_255;
assign enable_check_to_variable_255[0] = enable_check_95_to_variable_255;
// 将变量节点255的输出与校验节点95的输入相连
assign value_variable_255_to_check_95 = value_variable_255_to_check[5:0];
assign enable_variable_255_to_check_95 = enable_variable_255_to_check;

// 对校验节点111传递过来的数据进行整合
assign value_check_to_variable_255[11:6] = value_check_111_to_variable_255;
assign enable_check_to_variable_255[1] = enable_check_111_to_variable_255;
// 将变量节点255的输出与校验节点111的输入相连
assign value_variable_255_to_check_111 = value_variable_255_to_check[11:6];
assign enable_variable_255_to_check_111 = enable_variable_255_to_check;

// 对校验节点122传递过来的数据进行整合
assign value_check_to_variable_255[17:12] = value_check_122_to_variable_255;
assign enable_check_to_variable_255[2] = enable_check_122_to_variable_255;
// 将变量节点255的输出与校验节点122的输入相连
assign value_variable_255_to_check_122 = value_variable_255_to_check[17:12];
assign enable_variable_255_to_check_122 = enable_variable_255_to_check;


// 校验节点0
Check_Node #(.weight(6),.length(6)) u_Check_Node_0(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_0),
.variable_enable_input(enable_check_to_variable_0),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_0_to_check),
.check_enable_output(enable_variable_0_to_check)
);

// 校验节点1
Check_Node #(.weight(6),.length(6)) u_Check_Node_1(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_1),
.variable_enable_input(enable_check_to_variable_1),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_1_to_check),
.check_enable_output(enable_variable_1_to_check)
);

// 校验节点2
Check_Node #(.weight(6),.length(6)) u_Check_Node_2(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_2),
.variable_enable_input(enable_check_to_variable_2),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_2_to_check),
.check_enable_output(enable_variable_2_to_check)
);

// 校验节点3
Check_Node #(.weight(6),.length(6)) u_Check_Node_3(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_3),
.variable_enable_input(enable_check_to_variable_3),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_3_to_check),
.check_enable_output(enable_variable_3_to_check)
);

// 校验节点4
Check_Node #(.weight(6),.length(6)) u_Check_Node_4(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_4),
.variable_enable_input(enable_check_to_variable_4),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_4_to_check),
.check_enable_output(enable_variable_4_to_check)
);

// 校验节点5
Check_Node #(.weight(6),.length(6)) u_Check_Node_5(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_5),
.variable_enable_input(enable_check_to_variable_5),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_5_to_check),
.check_enable_output(enable_variable_5_to_check)
);

// 校验节点6
Check_Node #(.weight(6),.length(6)) u_Check_Node_6(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_6),
.variable_enable_input(enable_check_to_variable_6),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_6_to_check),
.check_enable_output(enable_variable_6_to_check)
);

// 校验节点7
Check_Node #(.weight(6),.length(6)) u_Check_Node_7(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_7),
.variable_enable_input(enable_check_to_variable_7),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_7_to_check),
.check_enable_output(enable_variable_7_to_check)
);

// 校验节点8
Check_Node #(.weight(6),.length(6)) u_Check_Node_8(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_8),
.variable_enable_input(enable_check_to_variable_8),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_8_to_check),
.check_enable_output(enable_variable_8_to_check)
);

// 校验节点9
Check_Node #(.weight(6),.length(6)) u_Check_Node_9(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_9),
.variable_enable_input(enable_check_to_variable_9),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_9_to_check),
.check_enable_output(enable_variable_9_to_check)
);

// 校验节点10
Check_Node #(.weight(6),.length(6)) u_Check_Node_10(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_10),
.variable_enable_input(enable_check_to_variable_10),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_10_to_check),
.check_enable_output(enable_variable_10_to_check)
);

// 校验节点11
Check_Node #(.weight(6),.length(6)) u_Check_Node_11(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_11),
.variable_enable_input(enable_check_to_variable_11),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_11_to_check),
.check_enable_output(enable_variable_11_to_check)
);

// 校验节点12
Check_Node #(.weight(6),.length(6)) u_Check_Node_12(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_12),
.variable_enable_input(enable_check_to_variable_12),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_12_to_check),
.check_enable_output(enable_variable_12_to_check)
);

// 校验节点13
Check_Node #(.weight(6),.length(6)) u_Check_Node_13(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_13),
.variable_enable_input(enable_check_to_variable_13),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_13_to_check),
.check_enable_output(enable_variable_13_to_check)
);

// 校验节点14
Check_Node #(.weight(6),.length(6)) u_Check_Node_14(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_14),
.variable_enable_input(enable_check_to_variable_14),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_14_to_check),
.check_enable_output(enable_variable_14_to_check)
);

// 校验节点15
Check_Node #(.weight(6),.length(6)) u_Check_Node_15(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_15),
.variable_enable_input(enable_check_to_variable_15),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_15_to_check),
.check_enable_output(enable_variable_15_to_check)
);

// 校验节点16
Check_Node #(.weight(6),.length(6)) u_Check_Node_16(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_16),
.variable_enable_input(enable_check_to_variable_16),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_16_to_check),
.check_enable_output(enable_variable_16_to_check)
);

// 校验节点17
Check_Node #(.weight(6),.length(6)) u_Check_Node_17(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_17),
.variable_enable_input(enable_check_to_variable_17),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_17_to_check),
.check_enable_output(enable_variable_17_to_check)
);

// 校验节点18
Check_Node #(.weight(6),.length(6)) u_Check_Node_18(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_18),
.variable_enable_input(enable_check_to_variable_18),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_18_to_check),
.check_enable_output(enable_variable_18_to_check)
);

// 校验节点19
Check_Node #(.weight(6),.length(6)) u_Check_Node_19(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_19),
.variable_enable_input(enable_check_to_variable_19),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_19_to_check),
.check_enable_output(enable_variable_19_to_check)
);

// 校验节点20
Check_Node #(.weight(6),.length(6)) u_Check_Node_20(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_20),
.variable_enable_input(enable_check_to_variable_20),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_20_to_check),
.check_enable_output(enable_variable_20_to_check)
);

// 校验节点21
Check_Node #(.weight(6),.length(6)) u_Check_Node_21(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_21),
.variable_enable_input(enable_check_to_variable_21),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_21_to_check),
.check_enable_output(enable_variable_21_to_check)
);

// 校验节点22
Check_Node #(.weight(6),.length(6)) u_Check_Node_22(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_22),
.variable_enable_input(enable_check_to_variable_22),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_22_to_check),
.check_enable_output(enable_variable_22_to_check)
);

// 校验节点23
Check_Node #(.weight(6),.length(6)) u_Check_Node_23(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_23),
.variable_enable_input(enable_check_to_variable_23),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_23_to_check),
.check_enable_output(enable_variable_23_to_check)
);

// 校验节点24
Check_Node #(.weight(6),.length(6)) u_Check_Node_24(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_24),
.variable_enable_input(enable_check_to_variable_24),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_24_to_check),
.check_enable_output(enable_variable_24_to_check)
);

// 校验节点25
Check_Node #(.weight(6),.length(6)) u_Check_Node_25(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_25),
.variable_enable_input(enable_check_to_variable_25),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_25_to_check),
.check_enable_output(enable_variable_25_to_check)
);

// 校验节点26
Check_Node #(.weight(6),.length(6)) u_Check_Node_26(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_26),
.variable_enable_input(enable_check_to_variable_26),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_26_to_check),
.check_enable_output(enable_variable_26_to_check)
);

// 校验节点27
Check_Node #(.weight(6),.length(6)) u_Check_Node_27(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_27),
.variable_enable_input(enable_check_to_variable_27),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_27_to_check),
.check_enable_output(enable_variable_27_to_check)
);

// 校验节点28
Check_Node #(.weight(6),.length(6)) u_Check_Node_28(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_28),
.variable_enable_input(enable_check_to_variable_28),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_28_to_check),
.check_enable_output(enable_variable_28_to_check)
);

// 校验节点29
Check_Node #(.weight(6),.length(6)) u_Check_Node_29(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_29),
.variable_enable_input(enable_check_to_variable_29),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_29_to_check),
.check_enable_output(enable_variable_29_to_check)
);

// 校验节点30
Check_Node #(.weight(6),.length(6)) u_Check_Node_30(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_30),
.variable_enable_input(enable_check_to_variable_30),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_30_to_check),
.check_enable_output(enable_variable_30_to_check)
);

// 校验节点31
Check_Node #(.weight(6),.length(6)) u_Check_Node_31(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_31),
.variable_enable_input(enable_check_to_variable_31),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_31_to_check),
.check_enable_output(enable_variable_31_to_check)
);

// 校验节点32
Check_Node #(.weight(6),.length(6)) u_Check_Node_32(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_32),
.variable_enable_input(enable_check_to_variable_32),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_32_to_check),
.check_enable_output(enable_variable_32_to_check)
);

// 校验节点33
Check_Node #(.weight(6),.length(6)) u_Check_Node_33(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_33),
.variable_enable_input(enable_check_to_variable_33),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_33_to_check),
.check_enable_output(enable_variable_33_to_check)
);

// 校验节点34
Check_Node #(.weight(6),.length(6)) u_Check_Node_34(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_34),
.variable_enable_input(enable_check_to_variable_34),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_34_to_check),
.check_enable_output(enable_variable_34_to_check)
);

// 校验节点35
Check_Node #(.weight(6),.length(6)) u_Check_Node_35(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_35),
.variable_enable_input(enable_check_to_variable_35),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_35_to_check),
.check_enable_output(enable_variable_35_to_check)
);

// 校验节点36
Check_Node #(.weight(6),.length(6)) u_Check_Node_36(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_36),
.variable_enable_input(enable_check_to_variable_36),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_36_to_check),
.check_enable_output(enable_variable_36_to_check)
);

// 校验节点37
Check_Node #(.weight(6),.length(6)) u_Check_Node_37(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_37),
.variable_enable_input(enable_check_to_variable_37),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_37_to_check),
.check_enable_output(enable_variable_37_to_check)
);

// 校验节点38
Check_Node #(.weight(6),.length(6)) u_Check_Node_38(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_38),
.variable_enable_input(enable_check_to_variable_38),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_38_to_check),
.check_enable_output(enable_variable_38_to_check)
);

// 校验节点39
Check_Node #(.weight(6),.length(6)) u_Check_Node_39(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_39),
.variable_enable_input(enable_check_to_variable_39),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_39_to_check),
.check_enable_output(enable_variable_39_to_check)
);

// 校验节点40
Check_Node #(.weight(6),.length(6)) u_Check_Node_40(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_40),
.variable_enable_input(enable_check_to_variable_40),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_40_to_check),
.check_enable_output(enable_variable_40_to_check)
);

// 校验节点41
Check_Node #(.weight(6),.length(6)) u_Check_Node_41(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_41),
.variable_enable_input(enable_check_to_variable_41),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_41_to_check),
.check_enable_output(enable_variable_41_to_check)
);

// 校验节点42
Check_Node #(.weight(6),.length(6)) u_Check_Node_42(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_42),
.variable_enable_input(enable_check_to_variable_42),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_42_to_check),
.check_enable_output(enable_variable_42_to_check)
);

// 校验节点43
Check_Node #(.weight(6),.length(6)) u_Check_Node_43(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_43),
.variable_enable_input(enable_check_to_variable_43),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_43_to_check),
.check_enable_output(enable_variable_43_to_check)
);

// 校验节点44
Check_Node #(.weight(6),.length(6)) u_Check_Node_44(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_44),
.variable_enable_input(enable_check_to_variable_44),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_44_to_check),
.check_enable_output(enable_variable_44_to_check)
);

// 校验节点45
Check_Node #(.weight(6),.length(6)) u_Check_Node_45(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_45),
.variable_enable_input(enable_check_to_variable_45),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_45_to_check),
.check_enable_output(enable_variable_45_to_check)
);

// 校验节点46
Check_Node #(.weight(6),.length(6)) u_Check_Node_46(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_46),
.variable_enable_input(enable_check_to_variable_46),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_46_to_check),
.check_enable_output(enable_variable_46_to_check)
);

// 校验节点47
Check_Node #(.weight(6),.length(6)) u_Check_Node_47(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_47),
.variable_enable_input(enable_check_to_variable_47),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_47_to_check),
.check_enable_output(enable_variable_47_to_check)
);

// 校验节点48
Check_Node #(.weight(6),.length(6)) u_Check_Node_48(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_48),
.variable_enable_input(enable_check_to_variable_48),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_48_to_check),
.check_enable_output(enable_variable_48_to_check)
);

// 校验节点49
Check_Node #(.weight(6),.length(6)) u_Check_Node_49(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_49),
.variable_enable_input(enable_check_to_variable_49),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_49_to_check),
.check_enable_output(enable_variable_49_to_check)
);

// 校验节点50
Check_Node #(.weight(6),.length(6)) u_Check_Node_50(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_50),
.variable_enable_input(enable_check_to_variable_50),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_50_to_check),
.check_enable_output(enable_variable_50_to_check)
);

// 校验节点51
Check_Node #(.weight(6),.length(6)) u_Check_Node_51(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_51),
.variable_enable_input(enable_check_to_variable_51),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_51_to_check),
.check_enable_output(enable_variable_51_to_check)
);

// 校验节点52
Check_Node #(.weight(6),.length(6)) u_Check_Node_52(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_52),
.variable_enable_input(enable_check_to_variable_52),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_52_to_check),
.check_enable_output(enable_variable_52_to_check)
);

// 校验节点53
Check_Node #(.weight(6),.length(6)) u_Check_Node_53(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_53),
.variable_enable_input(enable_check_to_variable_53),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_53_to_check),
.check_enable_output(enable_variable_53_to_check)
);

// 校验节点54
Check_Node #(.weight(6),.length(6)) u_Check_Node_54(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_54),
.variable_enable_input(enable_check_to_variable_54),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_54_to_check),
.check_enable_output(enable_variable_54_to_check)
);

// 校验节点55
Check_Node #(.weight(6),.length(6)) u_Check_Node_55(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_55),
.variable_enable_input(enable_check_to_variable_55),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_55_to_check),
.check_enable_output(enable_variable_55_to_check)
);

// 校验节点56
Check_Node #(.weight(6),.length(6)) u_Check_Node_56(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_56),
.variable_enable_input(enable_check_to_variable_56),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_56_to_check),
.check_enable_output(enable_variable_56_to_check)
);

// 校验节点57
Check_Node #(.weight(6),.length(6)) u_Check_Node_57(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_57),
.variable_enable_input(enable_check_to_variable_57),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_57_to_check),
.check_enable_output(enable_variable_57_to_check)
);

// 校验节点58
Check_Node #(.weight(6),.length(6)) u_Check_Node_58(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_58),
.variable_enable_input(enable_check_to_variable_58),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_58_to_check),
.check_enable_output(enable_variable_58_to_check)
);

// 校验节点59
Check_Node #(.weight(6),.length(6)) u_Check_Node_59(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_59),
.variable_enable_input(enable_check_to_variable_59),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_59_to_check),
.check_enable_output(enable_variable_59_to_check)
);

// 校验节点60
Check_Node #(.weight(6),.length(6)) u_Check_Node_60(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_60),
.variable_enable_input(enable_check_to_variable_60),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_60_to_check),
.check_enable_output(enable_variable_60_to_check)
);

// 校验节点61
Check_Node #(.weight(6),.length(6)) u_Check_Node_61(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_61),
.variable_enable_input(enable_check_to_variable_61),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_61_to_check),
.check_enable_output(enable_variable_61_to_check)
);

// 校验节点62
Check_Node #(.weight(6),.length(6)) u_Check_Node_62(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_62),
.variable_enable_input(enable_check_to_variable_62),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_62_to_check),
.check_enable_output(enable_variable_62_to_check)
);

// 校验节点63
Check_Node #(.weight(6),.length(6)) u_Check_Node_63(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_63),
.variable_enable_input(enable_check_to_variable_63),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_63_to_check),
.check_enable_output(enable_variable_63_to_check)
);

// 校验节点64
Check_Node #(.weight(6),.length(6)) u_Check_Node_64(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_64),
.variable_enable_input(enable_check_to_variable_64),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_64_to_check),
.check_enable_output(enable_variable_64_to_check)
);

// 校验节点65
Check_Node #(.weight(6),.length(6)) u_Check_Node_65(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_65),
.variable_enable_input(enable_check_to_variable_65),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_65_to_check),
.check_enable_output(enable_variable_65_to_check)
);

// 校验节点66
Check_Node #(.weight(6),.length(6)) u_Check_Node_66(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_66),
.variable_enable_input(enable_check_to_variable_66),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_66_to_check),
.check_enable_output(enable_variable_66_to_check)
);

// 校验节点67
Check_Node #(.weight(6),.length(6)) u_Check_Node_67(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_67),
.variable_enable_input(enable_check_to_variable_67),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_67_to_check),
.check_enable_output(enable_variable_67_to_check)
);

// 校验节点68
Check_Node #(.weight(6),.length(6)) u_Check_Node_68(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_68),
.variable_enable_input(enable_check_to_variable_68),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_68_to_check),
.check_enable_output(enable_variable_68_to_check)
);

// 校验节点69
Check_Node #(.weight(6),.length(6)) u_Check_Node_69(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_69),
.variable_enable_input(enable_check_to_variable_69),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_69_to_check),
.check_enable_output(enable_variable_69_to_check)
);

// 校验节点70
Check_Node #(.weight(6),.length(6)) u_Check_Node_70(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_70),
.variable_enable_input(enable_check_to_variable_70),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_70_to_check),
.check_enable_output(enable_variable_70_to_check)
);

// 校验节点71
Check_Node #(.weight(6),.length(6)) u_Check_Node_71(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_71),
.variable_enable_input(enable_check_to_variable_71),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_71_to_check),
.check_enable_output(enable_variable_71_to_check)
);

// 校验节点72
Check_Node #(.weight(6),.length(6)) u_Check_Node_72(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_72),
.variable_enable_input(enable_check_to_variable_72),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_72_to_check),
.check_enable_output(enable_variable_72_to_check)
);

// 校验节点73
Check_Node #(.weight(6),.length(6)) u_Check_Node_73(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_73),
.variable_enable_input(enable_check_to_variable_73),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_73_to_check),
.check_enable_output(enable_variable_73_to_check)
);

// 校验节点74
Check_Node #(.weight(6),.length(6)) u_Check_Node_74(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_74),
.variable_enable_input(enable_check_to_variable_74),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_74_to_check),
.check_enable_output(enable_variable_74_to_check)
);

// 校验节点75
Check_Node #(.weight(6),.length(6)) u_Check_Node_75(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_75),
.variable_enable_input(enable_check_to_variable_75),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_75_to_check),
.check_enable_output(enable_variable_75_to_check)
);

// 校验节点76
Check_Node #(.weight(6),.length(6)) u_Check_Node_76(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_76),
.variable_enable_input(enable_check_to_variable_76),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_76_to_check),
.check_enable_output(enable_variable_76_to_check)
);

// 校验节点77
Check_Node #(.weight(6),.length(6)) u_Check_Node_77(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_77),
.variable_enable_input(enable_check_to_variable_77),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_77_to_check),
.check_enable_output(enable_variable_77_to_check)
);

// 校验节点78
Check_Node #(.weight(6),.length(6)) u_Check_Node_78(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_78),
.variable_enable_input(enable_check_to_variable_78),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_78_to_check),
.check_enable_output(enable_variable_78_to_check)
);

// 校验节点79
Check_Node #(.weight(6),.length(6)) u_Check_Node_79(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_79),
.variable_enable_input(enable_check_to_variable_79),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_79_to_check),
.check_enable_output(enable_variable_79_to_check)
);

// 校验节点80
Check_Node #(.weight(6),.length(6)) u_Check_Node_80(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_80),
.variable_enable_input(enable_check_to_variable_80),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_80_to_check),
.check_enable_output(enable_variable_80_to_check)
);

// 校验节点81
Check_Node #(.weight(6),.length(6)) u_Check_Node_81(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_81),
.variable_enable_input(enable_check_to_variable_81),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_81_to_check),
.check_enable_output(enable_variable_81_to_check)
);

// 校验节点82
Check_Node #(.weight(6),.length(6)) u_Check_Node_82(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_82),
.variable_enable_input(enable_check_to_variable_82),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_82_to_check),
.check_enable_output(enable_variable_82_to_check)
);

// 校验节点83
Check_Node #(.weight(6),.length(6)) u_Check_Node_83(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_83),
.variable_enable_input(enable_check_to_variable_83),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_83_to_check),
.check_enable_output(enable_variable_83_to_check)
);

// 校验节点84
Check_Node #(.weight(6),.length(6)) u_Check_Node_84(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_84),
.variable_enable_input(enable_check_to_variable_84),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_84_to_check),
.check_enable_output(enable_variable_84_to_check)
);

// 校验节点85
Check_Node #(.weight(6),.length(6)) u_Check_Node_85(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_85),
.variable_enable_input(enable_check_to_variable_85),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_85_to_check),
.check_enable_output(enable_variable_85_to_check)
);

// 校验节点86
Check_Node #(.weight(6),.length(6)) u_Check_Node_86(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_86),
.variable_enable_input(enable_check_to_variable_86),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_86_to_check),
.check_enable_output(enable_variable_86_to_check)
);

// 校验节点87
Check_Node #(.weight(6),.length(6)) u_Check_Node_87(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_87),
.variable_enable_input(enable_check_to_variable_87),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_87_to_check),
.check_enable_output(enable_variable_87_to_check)
);

// 校验节点88
Check_Node #(.weight(6),.length(6)) u_Check_Node_88(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_88),
.variable_enable_input(enable_check_to_variable_88),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_88_to_check),
.check_enable_output(enable_variable_88_to_check)
);

// 校验节点89
Check_Node #(.weight(6),.length(6)) u_Check_Node_89(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_89),
.variable_enable_input(enable_check_to_variable_89),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_89_to_check),
.check_enable_output(enable_variable_89_to_check)
);

// 校验节点90
Check_Node #(.weight(6),.length(6)) u_Check_Node_90(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_90),
.variable_enable_input(enable_check_to_variable_90),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_90_to_check),
.check_enable_output(enable_variable_90_to_check)
);

// 校验节点91
Check_Node #(.weight(6),.length(6)) u_Check_Node_91(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_91),
.variable_enable_input(enable_check_to_variable_91),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_91_to_check),
.check_enable_output(enable_variable_91_to_check)
);

// 校验节点92
Check_Node #(.weight(6),.length(6)) u_Check_Node_92(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_92),
.variable_enable_input(enable_check_to_variable_92),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_92_to_check),
.check_enable_output(enable_variable_92_to_check)
);

// 校验节点93
Check_Node #(.weight(6),.length(6)) u_Check_Node_93(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_93),
.variable_enable_input(enable_check_to_variable_93),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_93_to_check),
.check_enable_output(enable_variable_93_to_check)
);

// 校验节点94
Check_Node #(.weight(6),.length(6)) u_Check_Node_94(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_94),
.variable_enable_input(enable_check_to_variable_94),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_94_to_check),
.check_enable_output(enable_variable_94_to_check)
);

// 校验节点95
Check_Node #(.weight(6),.length(6)) u_Check_Node_95(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_95),
.variable_enable_input(enable_check_to_variable_95),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_95_to_check),
.check_enable_output(enable_variable_95_to_check)
);

// 校验节点96
Check_Node #(.weight(6),.length(6)) u_Check_Node_96(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_96),
.variable_enable_input(enable_check_to_variable_96),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_96_to_check),
.check_enable_output(enable_variable_96_to_check)
);

// 校验节点97
Check_Node #(.weight(6),.length(6)) u_Check_Node_97(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_97),
.variable_enable_input(enable_check_to_variable_97),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_97_to_check),
.check_enable_output(enable_variable_97_to_check)
);

// 校验节点98
Check_Node #(.weight(6),.length(6)) u_Check_Node_98(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_98),
.variable_enable_input(enable_check_to_variable_98),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_98_to_check),
.check_enable_output(enable_variable_98_to_check)
);

// 校验节点99
Check_Node #(.weight(6),.length(6)) u_Check_Node_99(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_99),
.variable_enable_input(enable_check_to_variable_99),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_99_to_check),
.check_enable_output(enable_variable_99_to_check)
);

// 校验节点100
Check_Node #(.weight(6),.length(6)) u_Check_Node_100(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_100),
.variable_enable_input(enable_check_to_variable_100),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_100_to_check),
.check_enable_output(enable_variable_100_to_check)
);

// 校验节点101
Check_Node #(.weight(6),.length(6)) u_Check_Node_101(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_101),
.variable_enable_input(enable_check_to_variable_101),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_101_to_check),
.check_enable_output(enable_variable_101_to_check)
);

// 校验节点102
Check_Node #(.weight(6),.length(6)) u_Check_Node_102(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_102),
.variable_enable_input(enable_check_to_variable_102),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_102_to_check),
.check_enable_output(enable_variable_102_to_check)
);

// 校验节点103
Check_Node #(.weight(6),.length(6)) u_Check_Node_103(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_103),
.variable_enable_input(enable_check_to_variable_103),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_103_to_check),
.check_enable_output(enable_variable_103_to_check)
);

// 校验节点104
Check_Node #(.weight(6),.length(6)) u_Check_Node_104(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_104),
.variable_enable_input(enable_check_to_variable_104),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_104_to_check),
.check_enable_output(enable_variable_104_to_check)
);

// 校验节点105
Check_Node #(.weight(6),.length(6)) u_Check_Node_105(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_105),
.variable_enable_input(enable_check_to_variable_105),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_105_to_check),
.check_enable_output(enable_variable_105_to_check)
);

// 校验节点106
Check_Node #(.weight(6),.length(6)) u_Check_Node_106(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_106),
.variable_enable_input(enable_check_to_variable_106),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_106_to_check),
.check_enable_output(enable_variable_106_to_check)
);

// 校验节点107
Check_Node #(.weight(6),.length(6)) u_Check_Node_107(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_107),
.variable_enable_input(enable_check_to_variable_107),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_107_to_check),
.check_enable_output(enable_variable_107_to_check)
);

// 校验节点108
Check_Node #(.weight(6),.length(6)) u_Check_Node_108(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_108),
.variable_enable_input(enable_check_to_variable_108),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_108_to_check),
.check_enable_output(enable_variable_108_to_check)
);

// 校验节点109
Check_Node #(.weight(6),.length(6)) u_Check_Node_109(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_109),
.variable_enable_input(enable_check_to_variable_109),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_109_to_check),
.check_enable_output(enable_variable_109_to_check)
);

// 校验节点110
Check_Node #(.weight(6),.length(6)) u_Check_Node_110(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_110),
.variable_enable_input(enable_check_to_variable_110),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_110_to_check),
.check_enable_output(enable_variable_110_to_check)
);

// 校验节点111
Check_Node #(.weight(6),.length(6)) u_Check_Node_111(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_111),
.variable_enable_input(enable_check_to_variable_111),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_111_to_check),
.check_enable_output(enable_variable_111_to_check)
);

// 校验节点112
Check_Node #(.weight(6),.length(6)) u_Check_Node_112(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_112),
.variable_enable_input(enable_check_to_variable_112),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_112_to_check),
.check_enable_output(enable_variable_112_to_check)
);

// 校验节点113
Check_Node #(.weight(6),.length(6)) u_Check_Node_113(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_113),
.variable_enable_input(enable_check_to_variable_113),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_113_to_check),
.check_enable_output(enable_variable_113_to_check)
);

// 校验节点114
Check_Node #(.weight(6),.length(6)) u_Check_Node_114(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_114),
.variable_enable_input(enable_check_to_variable_114),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_114_to_check),
.check_enable_output(enable_variable_114_to_check)
);

// 校验节点115
Check_Node #(.weight(6),.length(6)) u_Check_Node_115(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_115),
.variable_enable_input(enable_check_to_variable_115),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_115_to_check),
.check_enable_output(enable_variable_115_to_check)
);

// 校验节点116
Check_Node #(.weight(6),.length(6)) u_Check_Node_116(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_116),
.variable_enable_input(enable_check_to_variable_116),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_116_to_check),
.check_enable_output(enable_variable_116_to_check)
);

// 校验节点117
Check_Node #(.weight(6),.length(6)) u_Check_Node_117(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_117),
.variable_enable_input(enable_check_to_variable_117),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_117_to_check),
.check_enable_output(enable_variable_117_to_check)
);

// 校验节点118
Check_Node #(.weight(6),.length(6)) u_Check_Node_118(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_118),
.variable_enable_input(enable_check_to_variable_118),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_118_to_check),
.check_enable_output(enable_variable_118_to_check)
);

// 校验节点119
Check_Node #(.weight(6),.length(6)) u_Check_Node_119(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_119),
.variable_enable_input(enable_check_to_variable_119),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_119_to_check),
.check_enable_output(enable_variable_119_to_check)
);

// 校验节点120
Check_Node #(.weight(6),.length(6)) u_Check_Node_120(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_120),
.variable_enable_input(enable_check_to_variable_120),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_120_to_check),
.check_enable_output(enable_variable_120_to_check)
);

// 校验节点121
Check_Node #(.weight(6),.length(6)) u_Check_Node_121(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_121),
.variable_enable_input(enable_check_to_variable_121),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_121_to_check),
.check_enable_output(enable_variable_121_to_check)
);

// 校验节点122
Check_Node #(.weight(6),.length(6)) u_Check_Node_122(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_122),
.variable_enable_input(enable_check_to_variable_122),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_122_to_check),
.check_enable_output(enable_variable_122_to_check)
);

// 校验节点123
Check_Node #(.weight(6),.length(6)) u_Check_Node_123(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_123),
.variable_enable_input(enable_check_to_variable_123),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_123_to_check),
.check_enable_output(enable_variable_123_to_check)
);

// 校验节点124
Check_Node #(.weight(6),.length(6)) u_Check_Node_124(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_124),
.variable_enable_input(enable_check_to_variable_124),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_124_to_check),
.check_enable_output(enable_variable_124_to_check)
);

// 校验节点125
Check_Node #(.weight(6),.length(6)) u_Check_Node_125(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_125),
.variable_enable_input(enable_check_to_variable_125),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_125_to_check),
.check_enable_output(enable_variable_125_to_check)
);

// 校验节点126
Check_Node #(.weight(6),.length(6)) u_Check_Node_126(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_126),
.variable_enable_input(enable_check_to_variable_126),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_126_to_check),
.check_enable_output(enable_variable_126_to_check)
);

// 校验节点127
Check_Node #(.weight(6),.length(6)) u_Check_Node_127(
.clk(clk),
.rst(rst),
.check_begin(check_begin),
.variable_value_input(value_check_to_variable_127),
.variable_enable_input(enable_check_to_variable_127),
.decision_down(),
.decision_success(),
.decision_down_receive(),
.check_value_output(value_variable_127_to_check),
.check_enable_output(enable_variable_127_to_check)
);


// 变量节点0
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_0(
.clk(clk),
.rst(rst),
.initial_value(initial_value[0]),
.initial_value_enable(initial_value_enable[0]),
.initial_down(initial_down[0]),
.check_value_input(value_check_to_variable_0),
.check_enable_input(enable_check_to_variable_0),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_0_to_decision),
.value_variable_to_check(value_variable_0_to_check),
.variable_enable(enable_variable_0_to_check)
);

// 变量节点1
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_1(
.clk(clk),
.rst(rst),
.initial_value(initial_value[1]),
.initial_value_enable(initial_value_enable[1]),
.initial_down(initial_down[1]),
.check_value_input(value_check_to_variable_1),
.check_enable_input(enable_check_to_variable_1),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_1_to_decision),
.value_variable_to_check(value_variable_1_to_check),
.variable_enable(enable_variable_1_to_check)
);

// 变量节点2
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_2(
.clk(clk),
.rst(rst),
.initial_value(initial_value[2]),
.initial_value_enable(initial_value_enable[2]),
.initial_down(initial_down[2]),
.check_value_input(value_check_to_variable_2),
.check_enable_input(enable_check_to_variable_2),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_2_to_decision),
.value_variable_to_check(value_variable_2_to_check),
.variable_enable(enable_variable_2_to_check)
);

// 变量节点3
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_3(
.clk(clk),
.rst(rst),
.initial_value(initial_value[3]),
.initial_value_enable(initial_value_enable[3]),
.initial_down(initial_down[3]),
.check_value_input(value_check_to_variable_3),
.check_enable_input(enable_check_to_variable_3),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_3_to_decision),
.value_variable_to_check(value_variable_3_to_check),
.variable_enable(enable_variable_3_to_check)
);

// 变量节点4
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_4(
.clk(clk),
.rst(rst),
.initial_value(initial_value[4]),
.initial_value_enable(initial_value_enable[4]),
.initial_down(initial_down[4]),
.check_value_input(value_check_to_variable_4),
.check_enable_input(enable_check_to_variable_4),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_4_to_decision),
.value_variable_to_check(value_variable_4_to_check),
.variable_enable(enable_variable_4_to_check)
);

// 变量节点5
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_5(
.clk(clk),
.rst(rst),
.initial_value(initial_value[5]),
.initial_value_enable(initial_value_enable[5]),
.initial_down(initial_down[5]),
.check_value_input(value_check_to_variable_5),
.check_enable_input(enable_check_to_variable_5),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_5_to_decision),
.value_variable_to_check(value_variable_5_to_check),
.variable_enable(enable_variable_5_to_check)
);

// 变量节点6
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_6(
.clk(clk),
.rst(rst),
.initial_value(initial_value[6]),
.initial_value_enable(initial_value_enable[6]),
.initial_down(initial_down[6]),
.check_value_input(value_check_to_variable_6),
.check_enable_input(enable_check_to_variable_6),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_6_to_decision),
.value_variable_to_check(value_variable_6_to_check),
.variable_enable(enable_variable_6_to_check)
);

// 变量节点7
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_7(
.clk(clk),
.rst(rst),
.initial_value(initial_value[7]),
.initial_value_enable(initial_value_enable[7]),
.initial_down(initial_down[7]),
.check_value_input(value_check_to_variable_7),
.check_enable_input(enable_check_to_variable_7),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_7_to_decision),
.value_variable_to_check(value_variable_7_to_check),
.variable_enable(enable_variable_7_to_check)
);

// 变量节点8
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_8(
.clk(clk),
.rst(rst),
.initial_value(initial_value[8]),
.initial_value_enable(initial_value_enable[8]),
.initial_down(initial_down[8]),
.check_value_input(value_check_to_variable_8),
.check_enable_input(enable_check_to_variable_8),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_8_to_decision),
.value_variable_to_check(value_variable_8_to_check),
.variable_enable(enable_variable_8_to_check)
);

// 变量节点9
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_9(
.clk(clk),
.rst(rst),
.initial_value(initial_value[9]),
.initial_value_enable(initial_value_enable[9]),
.initial_down(initial_down[9]),
.check_value_input(value_check_to_variable_9),
.check_enable_input(enable_check_to_variable_9),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_9_to_decision),
.value_variable_to_check(value_variable_9_to_check),
.variable_enable(enable_variable_9_to_check)
);

// 变量节点10
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_10(
.clk(clk),
.rst(rst),
.initial_value(initial_value[10]),
.initial_value_enable(initial_value_enable[10]),
.initial_down(initial_down[10]),
.check_value_input(value_check_to_variable_10),
.check_enable_input(enable_check_to_variable_10),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_10_to_decision),
.value_variable_to_check(value_variable_10_to_check),
.variable_enable(enable_variable_10_to_check)
);

// 变量节点11
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_11(
.clk(clk),
.rst(rst),
.initial_value(initial_value[11]),
.initial_value_enable(initial_value_enable[11]),
.initial_down(initial_down[11]),
.check_value_input(value_check_to_variable_11),
.check_enable_input(enable_check_to_variable_11),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_11_to_decision),
.value_variable_to_check(value_variable_11_to_check),
.variable_enable(enable_variable_11_to_check)
);

// 变量节点12
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_12(
.clk(clk),
.rst(rst),
.initial_value(initial_value[12]),
.initial_value_enable(initial_value_enable[12]),
.initial_down(initial_down[12]),
.check_value_input(value_check_to_variable_12),
.check_enable_input(enable_check_to_variable_12),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_12_to_decision),
.value_variable_to_check(value_variable_12_to_check),
.variable_enable(enable_variable_12_to_check)
);

// 变量节点13
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_13(
.clk(clk),
.rst(rst),
.initial_value(initial_value[13]),
.initial_value_enable(initial_value_enable[13]),
.initial_down(initial_down[13]),
.check_value_input(value_check_to_variable_13),
.check_enable_input(enable_check_to_variable_13),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_13_to_decision),
.value_variable_to_check(value_variable_13_to_check),
.variable_enable(enable_variable_13_to_check)
);

// 变量节点14
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_14(
.clk(clk),
.rst(rst),
.initial_value(initial_value[14]),
.initial_value_enable(initial_value_enable[14]),
.initial_down(initial_down[14]),
.check_value_input(value_check_to_variable_14),
.check_enable_input(enable_check_to_variable_14),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_14_to_decision),
.value_variable_to_check(value_variable_14_to_check),
.variable_enable(enable_variable_14_to_check)
);

// 变量节点15
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_15(
.clk(clk),
.rst(rst),
.initial_value(initial_value[15]),
.initial_value_enable(initial_value_enable[15]),
.initial_down(initial_down[15]),
.check_value_input(value_check_to_variable_15),
.check_enable_input(enable_check_to_variable_15),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_15_to_decision),
.value_variable_to_check(value_variable_15_to_check),
.variable_enable(enable_variable_15_to_check)
);

// 变量节点16
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_16(
.clk(clk),
.rst(rst),
.initial_value(initial_value[16]),
.initial_value_enable(initial_value_enable[16]),
.initial_down(initial_down[16]),
.check_value_input(value_check_to_variable_16),
.check_enable_input(enable_check_to_variable_16),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_16_to_decision),
.value_variable_to_check(value_variable_16_to_check),
.variable_enable(enable_variable_16_to_check)
);

// 变量节点17
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_17(
.clk(clk),
.rst(rst),
.initial_value(initial_value[17]),
.initial_value_enable(initial_value_enable[17]),
.initial_down(initial_down[17]),
.check_value_input(value_check_to_variable_17),
.check_enable_input(enable_check_to_variable_17),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_17_to_decision),
.value_variable_to_check(value_variable_17_to_check),
.variable_enable(enable_variable_17_to_check)
);

// 变量节点18
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_18(
.clk(clk),
.rst(rst),
.initial_value(initial_value[18]),
.initial_value_enable(initial_value_enable[18]),
.initial_down(initial_down[18]),
.check_value_input(value_check_to_variable_18),
.check_enable_input(enable_check_to_variable_18),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_18_to_decision),
.value_variable_to_check(value_variable_18_to_check),
.variable_enable(enable_variable_18_to_check)
);

// 变量节点19
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_19(
.clk(clk),
.rst(rst),
.initial_value(initial_value[19]),
.initial_value_enable(initial_value_enable[19]),
.initial_down(initial_down[19]),
.check_value_input(value_check_to_variable_19),
.check_enable_input(enable_check_to_variable_19),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_19_to_decision),
.value_variable_to_check(value_variable_19_to_check),
.variable_enable(enable_variable_19_to_check)
);

// 变量节点20
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_20(
.clk(clk),
.rst(rst),
.initial_value(initial_value[20]),
.initial_value_enable(initial_value_enable[20]),
.initial_down(initial_down[20]),
.check_value_input(value_check_to_variable_20),
.check_enable_input(enable_check_to_variable_20),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_20_to_decision),
.value_variable_to_check(value_variable_20_to_check),
.variable_enable(enable_variable_20_to_check)
);

// 变量节点21
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_21(
.clk(clk),
.rst(rst),
.initial_value(initial_value[21]),
.initial_value_enable(initial_value_enable[21]),
.initial_down(initial_down[21]),
.check_value_input(value_check_to_variable_21),
.check_enable_input(enable_check_to_variable_21),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_21_to_decision),
.value_variable_to_check(value_variable_21_to_check),
.variable_enable(enable_variable_21_to_check)
);

// 变量节点22
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_22(
.clk(clk),
.rst(rst),
.initial_value(initial_value[22]),
.initial_value_enable(initial_value_enable[22]),
.initial_down(initial_down[22]),
.check_value_input(value_check_to_variable_22),
.check_enable_input(enable_check_to_variable_22),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_22_to_decision),
.value_variable_to_check(value_variable_22_to_check),
.variable_enable(enable_variable_22_to_check)
);

// 变量节点23
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_23(
.clk(clk),
.rst(rst),
.initial_value(initial_value[23]),
.initial_value_enable(initial_value_enable[23]),
.initial_down(initial_down[23]),
.check_value_input(value_check_to_variable_23),
.check_enable_input(enable_check_to_variable_23),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_23_to_decision),
.value_variable_to_check(value_variable_23_to_check),
.variable_enable(enable_variable_23_to_check)
);

// 变量节点24
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_24(
.clk(clk),
.rst(rst),
.initial_value(initial_value[24]),
.initial_value_enable(initial_value_enable[24]),
.initial_down(initial_down[24]),
.check_value_input(value_check_to_variable_24),
.check_enable_input(enable_check_to_variable_24),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_24_to_decision),
.value_variable_to_check(value_variable_24_to_check),
.variable_enable(enable_variable_24_to_check)
);

// 变量节点25
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_25(
.clk(clk),
.rst(rst),
.initial_value(initial_value[25]),
.initial_value_enable(initial_value_enable[25]),
.initial_down(initial_down[25]),
.check_value_input(value_check_to_variable_25),
.check_enable_input(enable_check_to_variable_25),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_25_to_decision),
.value_variable_to_check(value_variable_25_to_check),
.variable_enable(enable_variable_25_to_check)
);

// 变量节点26
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_26(
.clk(clk),
.rst(rst),
.initial_value(initial_value[26]),
.initial_value_enable(initial_value_enable[26]),
.initial_down(initial_down[26]),
.check_value_input(value_check_to_variable_26),
.check_enable_input(enable_check_to_variable_26),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_26_to_decision),
.value_variable_to_check(value_variable_26_to_check),
.variable_enable(enable_variable_26_to_check)
);

// 变量节点27
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_27(
.clk(clk),
.rst(rst),
.initial_value(initial_value[27]),
.initial_value_enable(initial_value_enable[27]),
.initial_down(initial_down[27]),
.check_value_input(value_check_to_variable_27),
.check_enable_input(enable_check_to_variable_27),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_27_to_decision),
.value_variable_to_check(value_variable_27_to_check),
.variable_enable(enable_variable_27_to_check)
);

// 变量节点28
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_28(
.clk(clk),
.rst(rst),
.initial_value(initial_value[28]),
.initial_value_enable(initial_value_enable[28]),
.initial_down(initial_down[28]),
.check_value_input(value_check_to_variable_28),
.check_enable_input(enable_check_to_variable_28),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_28_to_decision),
.value_variable_to_check(value_variable_28_to_check),
.variable_enable(enable_variable_28_to_check)
);

// 变量节点29
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_29(
.clk(clk),
.rst(rst),
.initial_value(initial_value[29]),
.initial_value_enable(initial_value_enable[29]),
.initial_down(initial_down[29]),
.check_value_input(value_check_to_variable_29),
.check_enable_input(enable_check_to_variable_29),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_29_to_decision),
.value_variable_to_check(value_variable_29_to_check),
.variable_enable(enable_variable_29_to_check)
);

// 变量节点30
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_30(
.clk(clk),
.rst(rst),
.initial_value(initial_value[30]),
.initial_value_enable(initial_value_enable[30]),
.initial_down(initial_down[30]),
.check_value_input(value_check_to_variable_30),
.check_enable_input(enable_check_to_variable_30),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_30_to_decision),
.value_variable_to_check(value_variable_30_to_check),
.variable_enable(enable_variable_30_to_check)
);

// 变量节点31
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_31(
.clk(clk),
.rst(rst),
.initial_value(initial_value[31]),
.initial_value_enable(initial_value_enable[31]),
.initial_down(initial_down[31]),
.check_value_input(value_check_to_variable_31),
.check_enable_input(enable_check_to_variable_31),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_31_to_decision),
.value_variable_to_check(value_variable_31_to_check),
.variable_enable(enable_variable_31_to_check)
);

// 变量节点32
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_32(
.clk(clk),
.rst(rst),
.initial_value(initial_value[32]),
.initial_value_enable(initial_value_enable[32]),
.initial_down(initial_down[32]),
.check_value_input(value_check_to_variable_32),
.check_enable_input(enable_check_to_variable_32),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_32_to_decision),
.value_variable_to_check(value_variable_32_to_check),
.variable_enable(enable_variable_32_to_check)
);

// 变量节点33
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_33(
.clk(clk),
.rst(rst),
.initial_value(initial_value[33]),
.initial_value_enable(initial_value_enable[33]),
.initial_down(initial_down[33]),
.check_value_input(value_check_to_variable_33),
.check_enable_input(enable_check_to_variable_33),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_33_to_decision),
.value_variable_to_check(value_variable_33_to_check),
.variable_enable(enable_variable_33_to_check)
);

// 变量节点34
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_34(
.clk(clk),
.rst(rst),
.initial_value(initial_value[34]),
.initial_value_enable(initial_value_enable[34]),
.initial_down(initial_down[34]),
.check_value_input(value_check_to_variable_34),
.check_enable_input(enable_check_to_variable_34),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_34_to_decision),
.value_variable_to_check(value_variable_34_to_check),
.variable_enable(enable_variable_34_to_check)
);

// 变量节点35
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_35(
.clk(clk),
.rst(rst),
.initial_value(initial_value[35]),
.initial_value_enable(initial_value_enable[35]),
.initial_down(initial_down[35]),
.check_value_input(value_check_to_variable_35),
.check_enable_input(enable_check_to_variable_35),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_35_to_decision),
.value_variable_to_check(value_variable_35_to_check),
.variable_enable(enable_variable_35_to_check)
);

// 变量节点36
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_36(
.clk(clk),
.rst(rst),
.initial_value(initial_value[36]),
.initial_value_enable(initial_value_enable[36]),
.initial_down(initial_down[36]),
.check_value_input(value_check_to_variable_36),
.check_enable_input(enable_check_to_variable_36),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_36_to_decision),
.value_variable_to_check(value_variable_36_to_check),
.variable_enable(enable_variable_36_to_check)
);

// 变量节点37
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_37(
.clk(clk),
.rst(rst),
.initial_value(initial_value[37]),
.initial_value_enable(initial_value_enable[37]),
.initial_down(initial_down[37]),
.check_value_input(value_check_to_variable_37),
.check_enable_input(enable_check_to_variable_37),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_37_to_decision),
.value_variable_to_check(value_variable_37_to_check),
.variable_enable(enable_variable_37_to_check)
);

// 变量节点38
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_38(
.clk(clk),
.rst(rst),
.initial_value(initial_value[38]),
.initial_value_enable(initial_value_enable[38]),
.initial_down(initial_down[38]),
.check_value_input(value_check_to_variable_38),
.check_enable_input(enable_check_to_variable_38),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_38_to_decision),
.value_variable_to_check(value_variable_38_to_check),
.variable_enable(enable_variable_38_to_check)
);

// 变量节点39
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_39(
.clk(clk),
.rst(rst),
.initial_value(initial_value[39]),
.initial_value_enable(initial_value_enable[39]),
.initial_down(initial_down[39]),
.check_value_input(value_check_to_variable_39),
.check_enable_input(enable_check_to_variable_39),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_39_to_decision),
.value_variable_to_check(value_variable_39_to_check),
.variable_enable(enable_variable_39_to_check)
);

// 变量节点40
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_40(
.clk(clk),
.rst(rst),
.initial_value(initial_value[40]),
.initial_value_enable(initial_value_enable[40]),
.initial_down(initial_down[40]),
.check_value_input(value_check_to_variable_40),
.check_enable_input(enable_check_to_variable_40),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_40_to_decision),
.value_variable_to_check(value_variable_40_to_check),
.variable_enable(enable_variable_40_to_check)
);

// 变量节点41
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_41(
.clk(clk),
.rst(rst),
.initial_value(initial_value[41]),
.initial_value_enable(initial_value_enable[41]),
.initial_down(initial_down[41]),
.check_value_input(value_check_to_variable_41),
.check_enable_input(enable_check_to_variable_41),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_41_to_decision),
.value_variable_to_check(value_variable_41_to_check),
.variable_enable(enable_variable_41_to_check)
);

// 变量节点42
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_42(
.clk(clk),
.rst(rst),
.initial_value(initial_value[42]),
.initial_value_enable(initial_value_enable[42]),
.initial_down(initial_down[42]),
.check_value_input(value_check_to_variable_42),
.check_enable_input(enable_check_to_variable_42),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_42_to_decision),
.value_variable_to_check(value_variable_42_to_check),
.variable_enable(enable_variable_42_to_check)
);

// 变量节点43
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_43(
.clk(clk),
.rst(rst),
.initial_value(initial_value[43]),
.initial_value_enable(initial_value_enable[43]),
.initial_down(initial_down[43]),
.check_value_input(value_check_to_variable_43),
.check_enable_input(enable_check_to_variable_43),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_43_to_decision),
.value_variable_to_check(value_variable_43_to_check),
.variable_enable(enable_variable_43_to_check)
);

// 变量节点44
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_44(
.clk(clk),
.rst(rst),
.initial_value(initial_value[44]),
.initial_value_enable(initial_value_enable[44]),
.initial_down(initial_down[44]),
.check_value_input(value_check_to_variable_44),
.check_enable_input(enable_check_to_variable_44),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_44_to_decision),
.value_variable_to_check(value_variable_44_to_check),
.variable_enable(enable_variable_44_to_check)
);

// 变量节点45
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_45(
.clk(clk),
.rst(rst),
.initial_value(initial_value[45]),
.initial_value_enable(initial_value_enable[45]),
.initial_down(initial_down[45]),
.check_value_input(value_check_to_variable_45),
.check_enable_input(enable_check_to_variable_45),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_45_to_decision),
.value_variable_to_check(value_variable_45_to_check),
.variable_enable(enable_variable_45_to_check)
);

// 变量节点46
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_46(
.clk(clk),
.rst(rst),
.initial_value(initial_value[46]),
.initial_value_enable(initial_value_enable[46]),
.initial_down(initial_down[46]),
.check_value_input(value_check_to_variable_46),
.check_enable_input(enable_check_to_variable_46),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_46_to_decision),
.value_variable_to_check(value_variable_46_to_check),
.variable_enable(enable_variable_46_to_check)
);

// 变量节点47
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_47(
.clk(clk),
.rst(rst),
.initial_value(initial_value[47]),
.initial_value_enable(initial_value_enable[47]),
.initial_down(initial_down[47]),
.check_value_input(value_check_to_variable_47),
.check_enable_input(enable_check_to_variable_47),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_47_to_decision),
.value_variable_to_check(value_variable_47_to_check),
.variable_enable(enable_variable_47_to_check)
);

// 变量节点48
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_48(
.clk(clk),
.rst(rst),
.initial_value(initial_value[48]),
.initial_value_enable(initial_value_enable[48]),
.initial_down(initial_down[48]),
.check_value_input(value_check_to_variable_48),
.check_enable_input(enable_check_to_variable_48),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_48_to_decision),
.value_variable_to_check(value_variable_48_to_check),
.variable_enable(enable_variable_48_to_check)
);

// 变量节点49
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_49(
.clk(clk),
.rst(rst),
.initial_value(initial_value[49]),
.initial_value_enable(initial_value_enable[49]),
.initial_down(initial_down[49]),
.check_value_input(value_check_to_variable_49),
.check_enable_input(enable_check_to_variable_49),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_49_to_decision),
.value_variable_to_check(value_variable_49_to_check),
.variable_enable(enable_variable_49_to_check)
);

// 变量节点50
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_50(
.clk(clk),
.rst(rst),
.initial_value(initial_value[50]),
.initial_value_enable(initial_value_enable[50]),
.initial_down(initial_down[50]),
.check_value_input(value_check_to_variable_50),
.check_enable_input(enable_check_to_variable_50),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_50_to_decision),
.value_variable_to_check(value_variable_50_to_check),
.variable_enable(enable_variable_50_to_check)
);

// 变量节点51
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_51(
.clk(clk),
.rst(rst),
.initial_value(initial_value[51]),
.initial_value_enable(initial_value_enable[51]),
.initial_down(initial_down[51]),
.check_value_input(value_check_to_variable_51),
.check_enable_input(enable_check_to_variable_51),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_51_to_decision),
.value_variable_to_check(value_variable_51_to_check),
.variable_enable(enable_variable_51_to_check)
);

// 变量节点52
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_52(
.clk(clk),
.rst(rst),
.initial_value(initial_value[52]),
.initial_value_enable(initial_value_enable[52]),
.initial_down(initial_down[52]),
.check_value_input(value_check_to_variable_52),
.check_enable_input(enable_check_to_variable_52),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_52_to_decision),
.value_variable_to_check(value_variable_52_to_check),
.variable_enable(enable_variable_52_to_check)
);

// 变量节点53
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_53(
.clk(clk),
.rst(rst),
.initial_value(initial_value[53]),
.initial_value_enable(initial_value_enable[53]),
.initial_down(initial_down[53]),
.check_value_input(value_check_to_variable_53),
.check_enable_input(enable_check_to_variable_53),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_53_to_decision),
.value_variable_to_check(value_variable_53_to_check),
.variable_enable(enable_variable_53_to_check)
);

// 变量节点54
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_54(
.clk(clk),
.rst(rst),
.initial_value(initial_value[54]),
.initial_value_enable(initial_value_enable[54]),
.initial_down(initial_down[54]),
.check_value_input(value_check_to_variable_54),
.check_enable_input(enable_check_to_variable_54),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_54_to_decision),
.value_variable_to_check(value_variable_54_to_check),
.variable_enable(enable_variable_54_to_check)
);

// 变量节点55
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_55(
.clk(clk),
.rst(rst),
.initial_value(initial_value[55]),
.initial_value_enable(initial_value_enable[55]),
.initial_down(initial_down[55]),
.check_value_input(value_check_to_variable_55),
.check_enable_input(enable_check_to_variable_55),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_55_to_decision),
.value_variable_to_check(value_variable_55_to_check),
.variable_enable(enable_variable_55_to_check)
);

// 变量节点56
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_56(
.clk(clk),
.rst(rst),
.initial_value(initial_value[56]),
.initial_value_enable(initial_value_enable[56]),
.initial_down(initial_down[56]),
.check_value_input(value_check_to_variable_56),
.check_enable_input(enable_check_to_variable_56),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_56_to_decision),
.value_variable_to_check(value_variable_56_to_check),
.variable_enable(enable_variable_56_to_check)
);

// 变量节点57
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_57(
.clk(clk),
.rst(rst),
.initial_value(initial_value[57]),
.initial_value_enable(initial_value_enable[57]),
.initial_down(initial_down[57]),
.check_value_input(value_check_to_variable_57),
.check_enable_input(enable_check_to_variable_57),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_57_to_decision),
.value_variable_to_check(value_variable_57_to_check),
.variable_enable(enable_variable_57_to_check)
);

// 变量节点58
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_58(
.clk(clk),
.rst(rst),
.initial_value(initial_value[58]),
.initial_value_enable(initial_value_enable[58]),
.initial_down(initial_down[58]),
.check_value_input(value_check_to_variable_58),
.check_enable_input(enable_check_to_variable_58),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_58_to_decision),
.value_variable_to_check(value_variable_58_to_check),
.variable_enable(enable_variable_58_to_check)
);

// 变量节点59
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_59(
.clk(clk),
.rst(rst),
.initial_value(initial_value[59]),
.initial_value_enable(initial_value_enable[59]),
.initial_down(initial_down[59]),
.check_value_input(value_check_to_variable_59),
.check_enable_input(enable_check_to_variable_59),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_59_to_decision),
.value_variable_to_check(value_variable_59_to_check),
.variable_enable(enable_variable_59_to_check)
);

// 变量节点60
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_60(
.clk(clk),
.rst(rst),
.initial_value(initial_value[60]),
.initial_value_enable(initial_value_enable[60]),
.initial_down(initial_down[60]),
.check_value_input(value_check_to_variable_60),
.check_enable_input(enable_check_to_variable_60),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_60_to_decision),
.value_variable_to_check(value_variable_60_to_check),
.variable_enable(enable_variable_60_to_check)
);

// 变量节点61
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_61(
.clk(clk),
.rst(rst),
.initial_value(initial_value[61]),
.initial_value_enable(initial_value_enable[61]),
.initial_down(initial_down[61]),
.check_value_input(value_check_to_variable_61),
.check_enable_input(enable_check_to_variable_61),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_61_to_decision),
.value_variable_to_check(value_variable_61_to_check),
.variable_enable(enable_variable_61_to_check)
);

// 变量节点62
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_62(
.clk(clk),
.rst(rst),
.initial_value(initial_value[62]),
.initial_value_enable(initial_value_enable[62]),
.initial_down(initial_down[62]),
.check_value_input(value_check_to_variable_62),
.check_enable_input(enable_check_to_variable_62),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_62_to_decision),
.value_variable_to_check(value_variable_62_to_check),
.variable_enable(enable_variable_62_to_check)
);

// 变量节点63
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_63(
.clk(clk),
.rst(rst),
.initial_value(initial_value[63]),
.initial_value_enable(initial_value_enable[63]),
.initial_down(initial_down[63]),
.check_value_input(value_check_to_variable_63),
.check_enable_input(enable_check_to_variable_63),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_63_to_decision),
.value_variable_to_check(value_variable_63_to_check),
.variable_enable(enable_variable_63_to_check)
);

// 变量节点64
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_64(
.clk(clk),
.rst(rst),
.initial_value(initial_value[64]),
.initial_value_enable(initial_value_enable[64]),
.initial_down(initial_down[64]),
.check_value_input(value_check_to_variable_64),
.check_enable_input(enable_check_to_variable_64),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_64_to_decision),
.value_variable_to_check(value_variable_64_to_check),
.variable_enable(enable_variable_64_to_check)
);

// 变量节点65
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_65(
.clk(clk),
.rst(rst),
.initial_value(initial_value[65]),
.initial_value_enable(initial_value_enable[65]),
.initial_down(initial_down[65]),
.check_value_input(value_check_to_variable_65),
.check_enable_input(enable_check_to_variable_65),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_65_to_decision),
.value_variable_to_check(value_variable_65_to_check),
.variable_enable(enable_variable_65_to_check)
);

// 变量节点66
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_66(
.clk(clk),
.rst(rst),
.initial_value(initial_value[66]),
.initial_value_enable(initial_value_enable[66]),
.initial_down(initial_down[66]),
.check_value_input(value_check_to_variable_66),
.check_enable_input(enable_check_to_variable_66),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_66_to_decision),
.value_variable_to_check(value_variable_66_to_check),
.variable_enable(enable_variable_66_to_check)
);

// 变量节点67
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_67(
.clk(clk),
.rst(rst),
.initial_value(initial_value[67]),
.initial_value_enable(initial_value_enable[67]),
.initial_down(initial_down[67]),
.check_value_input(value_check_to_variable_67),
.check_enable_input(enable_check_to_variable_67),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_67_to_decision),
.value_variable_to_check(value_variable_67_to_check),
.variable_enable(enable_variable_67_to_check)
);

// 变量节点68
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_68(
.clk(clk),
.rst(rst),
.initial_value(initial_value[68]),
.initial_value_enable(initial_value_enable[68]),
.initial_down(initial_down[68]),
.check_value_input(value_check_to_variable_68),
.check_enable_input(enable_check_to_variable_68),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_68_to_decision),
.value_variable_to_check(value_variable_68_to_check),
.variable_enable(enable_variable_68_to_check)
);

// 变量节点69
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_69(
.clk(clk),
.rst(rst),
.initial_value(initial_value[69]),
.initial_value_enable(initial_value_enable[69]),
.initial_down(initial_down[69]),
.check_value_input(value_check_to_variable_69),
.check_enable_input(enable_check_to_variable_69),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_69_to_decision),
.value_variable_to_check(value_variable_69_to_check),
.variable_enable(enable_variable_69_to_check)
);

// 变量节点70
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_70(
.clk(clk),
.rst(rst),
.initial_value(initial_value[70]),
.initial_value_enable(initial_value_enable[70]),
.initial_down(initial_down[70]),
.check_value_input(value_check_to_variable_70),
.check_enable_input(enable_check_to_variable_70),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_70_to_decision),
.value_variable_to_check(value_variable_70_to_check),
.variable_enable(enable_variable_70_to_check)
);

// 变量节点71
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_71(
.clk(clk),
.rst(rst),
.initial_value(initial_value[71]),
.initial_value_enable(initial_value_enable[71]),
.initial_down(initial_down[71]),
.check_value_input(value_check_to_variable_71),
.check_enable_input(enable_check_to_variable_71),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_71_to_decision),
.value_variable_to_check(value_variable_71_to_check),
.variable_enable(enable_variable_71_to_check)
);

// 变量节点72
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_72(
.clk(clk),
.rst(rst),
.initial_value(initial_value[72]),
.initial_value_enable(initial_value_enable[72]),
.initial_down(initial_down[72]),
.check_value_input(value_check_to_variable_72),
.check_enable_input(enable_check_to_variable_72),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_72_to_decision),
.value_variable_to_check(value_variable_72_to_check),
.variable_enable(enable_variable_72_to_check)
);

// 变量节点73
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_73(
.clk(clk),
.rst(rst),
.initial_value(initial_value[73]),
.initial_value_enable(initial_value_enable[73]),
.initial_down(initial_down[73]),
.check_value_input(value_check_to_variable_73),
.check_enable_input(enable_check_to_variable_73),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_73_to_decision),
.value_variable_to_check(value_variable_73_to_check),
.variable_enable(enable_variable_73_to_check)
);

// 变量节点74
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_74(
.clk(clk),
.rst(rst),
.initial_value(initial_value[74]),
.initial_value_enable(initial_value_enable[74]),
.initial_down(initial_down[74]),
.check_value_input(value_check_to_variable_74),
.check_enable_input(enable_check_to_variable_74),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_74_to_decision),
.value_variable_to_check(value_variable_74_to_check),
.variable_enable(enable_variable_74_to_check)
);

// 变量节点75
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_75(
.clk(clk),
.rst(rst),
.initial_value(initial_value[75]),
.initial_value_enable(initial_value_enable[75]),
.initial_down(initial_down[75]),
.check_value_input(value_check_to_variable_75),
.check_enable_input(enable_check_to_variable_75),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_75_to_decision),
.value_variable_to_check(value_variable_75_to_check),
.variable_enable(enable_variable_75_to_check)
);

// 变量节点76
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_76(
.clk(clk),
.rst(rst),
.initial_value(initial_value[76]),
.initial_value_enable(initial_value_enable[76]),
.initial_down(initial_down[76]),
.check_value_input(value_check_to_variable_76),
.check_enable_input(enable_check_to_variable_76),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_76_to_decision),
.value_variable_to_check(value_variable_76_to_check),
.variable_enable(enable_variable_76_to_check)
);

// 变量节点77
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_77(
.clk(clk),
.rst(rst),
.initial_value(initial_value[77]),
.initial_value_enable(initial_value_enable[77]),
.initial_down(initial_down[77]),
.check_value_input(value_check_to_variable_77),
.check_enable_input(enable_check_to_variable_77),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_77_to_decision),
.value_variable_to_check(value_variable_77_to_check),
.variable_enable(enable_variable_77_to_check)
);

// 变量节点78
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_78(
.clk(clk),
.rst(rst),
.initial_value(initial_value[78]),
.initial_value_enable(initial_value_enable[78]),
.initial_down(initial_down[78]),
.check_value_input(value_check_to_variable_78),
.check_enable_input(enable_check_to_variable_78),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_78_to_decision),
.value_variable_to_check(value_variable_78_to_check),
.variable_enable(enable_variable_78_to_check)
);

// 变量节点79
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_79(
.clk(clk),
.rst(rst),
.initial_value(initial_value[79]),
.initial_value_enable(initial_value_enable[79]),
.initial_down(initial_down[79]),
.check_value_input(value_check_to_variable_79),
.check_enable_input(enable_check_to_variable_79),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_79_to_decision),
.value_variable_to_check(value_variable_79_to_check),
.variable_enable(enable_variable_79_to_check)
);

// 变量节点80
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_80(
.clk(clk),
.rst(rst),
.initial_value(initial_value[80]),
.initial_value_enable(initial_value_enable[80]),
.initial_down(initial_down[80]),
.check_value_input(value_check_to_variable_80),
.check_enable_input(enable_check_to_variable_80),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_80_to_decision),
.value_variable_to_check(value_variable_80_to_check),
.variable_enable(enable_variable_80_to_check)
);

// 变量节点81
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_81(
.clk(clk),
.rst(rst),
.initial_value(initial_value[81]),
.initial_value_enable(initial_value_enable[81]),
.initial_down(initial_down[81]),
.check_value_input(value_check_to_variable_81),
.check_enable_input(enable_check_to_variable_81),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_81_to_decision),
.value_variable_to_check(value_variable_81_to_check),
.variable_enable(enable_variable_81_to_check)
);

// 变量节点82
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_82(
.clk(clk),
.rst(rst),
.initial_value(initial_value[82]),
.initial_value_enable(initial_value_enable[82]),
.initial_down(initial_down[82]),
.check_value_input(value_check_to_variable_82),
.check_enable_input(enable_check_to_variable_82),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_82_to_decision),
.value_variable_to_check(value_variable_82_to_check),
.variable_enable(enable_variable_82_to_check)
);

// 变量节点83
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_83(
.clk(clk),
.rst(rst),
.initial_value(initial_value[83]),
.initial_value_enable(initial_value_enable[83]),
.initial_down(initial_down[83]),
.check_value_input(value_check_to_variable_83),
.check_enable_input(enable_check_to_variable_83),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_83_to_decision),
.value_variable_to_check(value_variable_83_to_check),
.variable_enable(enable_variable_83_to_check)
);

// 变量节点84
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_84(
.clk(clk),
.rst(rst),
.initial_value(initial_value[84]),
.initial_value_enable(initial_value_enable[84]),
.initial_down(initial_down[84]),
.check_value_input(value_check_to_variable_84),
.check_enable_input(enable_check_to_variable_84),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_84_to_decision),
.value_variable_to_check(value_variable_84_to_check),
.variable_enable(enable_variable_84_to_check)
);

// 变量节点85
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_85(
.clk(clk),
.rst(rst),
.initial_value(initial_value[85]),
.initial_value_enable(initial_value_enable[85]),
.initial_down(initial_down[85]),
.check_value_input(value_check_to_variable_85),
.check_enable_input(enable_check_to_variable_85),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_85_to_decision),
.value_variable_to_check(value_variable_85_to_check),
.variable_enable(enable_variable_85_to_check)
);

// 变量节点86
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_86(
.clk(clk),
.rst(rst),
.initial_value(initial_value[86]),
.initial_value_enable(initial_value_enable[86]),
.initial_down(initial_down[86]),
.check_value_input(value_check_to_variable_86),
.check_enable_input(enable_check_to_variable_86),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_86_to_decision),
.value_variable_to_check(value_variable_86_to_check),
.variable_enable(enable_variable_86_to_check)
);

// 变量节点87
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_87(
.clk(clk),
.rst(rst),
.initial_value(initial_value[87]),
.initial_value_enable(initial_value_enable[87]),
.initial_down(initial_down[87]),
.check_value_input(value_check_to_variable_87),
.check_enable_input(enable_check_to_variable_87),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_87_to_decision),
.value_variable_to_check(value_variable_87_to_check),
.variable_enable(enable_variable_87_to_check)
);

// 变量节点88
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_88(
.clk(clk),
.rst(rst),
.initial_value(initial_value[88]),
.initial_value_enable(initial_value_enable[88]),
.initial_down(initial_down[88]),
.check_value_input(value_check_to_variable_88),
.check_enable_input(enable_check_to_variable_88),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_88_to_decision),
.value_variable_to_check(value_variable_88_to_check),
.variable_enable(enable_variable_88_to_check)
);

// 变量节点89
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_89(
.clk(clk),
.rst(rst),
.initial_value(initial_value[89]),
.initial_value_enable(initial_value_enable[89]),
.initial_down(initial_down[89]),
.check_value_input(value_check_to_variable_89),
.check_enable_input(enable_check_to_variable_89),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_89_to_decision),
.value_variable_to_check(value_variable_89_to_check),
.variable_enable(enable_variable_89_to_check)
);

// 变量节点90
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_90(
.clk(clk),
.rst(rst),
.initial_value(initial_value[90]),
.initial_value_enable(initial_value_enable[90]),
.initial_down(initial_down[90]),
.check_value_input(value_check_to_variable_90),
.check_enable_input(enable_check_to_variable_90),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_90_to_decision),
.value_variable_to_check(value_variable_90_to_check),
.variable_enable(enable_variable_90_to_check)
);

// 变量节点91
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_91(
.clk(clk),
.rst(rst),
.initial_value(initial_value[91]),
.initial_value_enable(initial_value_enable[91]),
.initial_down(initial_down[91]),
.check_value_input(value_check_to_variable_91),
.check_enable_input(enable_check_to_variable_91),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_91_to_decision),
.value_variable_to_check(value_variable_91_to_check),
.variable_enable(enable_variable_91_to_check)
);

// 变量节点92
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_92(
.clk(clk),
.rst(rst),
.initial_value(initial_value[92]),
.initial_value_enable(initial_value_enable[92]),
.initial_down(initial_down[92]),
.check_value_input(value_check_to_variable_92),
.check_enable_input(enable_check_to_variable_92),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_92_to_decision),
.value_variable_to_check(value_variable_92_to_check),
.variable_enable(enable_variable_92_to_check)
);

// 变量节点93
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_93(
.clk(clk),
.rst(rst),
.initial_value(initial_value[93]),
.initial_value_enable(initial_value_enable[93]),
.initial_down(initial_down[93]),
.check_value_input(value_check_to_variable_93),
.check_enable_input(enable_check_to_variable_93),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_93_to_decision),
.value_variable_to_check(value_variable_93_to_check),
.variable_enable(enable_variable_93_to_check)
);

// 变量节点94
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_94(
.clk(clk),
.rst(rst),
.initial_value(initial_value[94]),
.initial_value_enable(initial_value_enable[94]),
.initial_down(initial_down[94]),
.check_value_input(value_check_to_variable_94),
.check_enable_input(enable_check_to_variable_94),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_94_to_decision),
.value_variable_to_check(value_variable_94_to_check),
.variable_enable(enable_variable_94_to_check)
);

// 变量节点95
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_95(
.clk(clk),
.rst(rst),
.initial_value(initial_value[95]),
.initial_value_enable(initial_value_enable[95]),
.initial_down(initial_down[95]),
.check_value_input(value_check_to_variable_95),
.check_enable_input(enable_check_to_variable_95),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_95_to_decision),
.value_variable_to_check(value_variable_95_to_check),
.variable_enable(enable_variable_95_to_check)
);

// 变量节点96
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_96(
.clk(clk),
.rst(rst),
.initial_value(initial_value[96]),
.initial_value_enable(initial_value_enable[96]),
.initial_down(initial_down[96]),
.check_value_input(value_check_to_variable_96),
.check_enable_input(enable_check_to_variable_96),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_96_to_decision),
.value_variable_to_check(value_variable_96_to_check),
.variable_enable(enable_variable_96_to_check)
);

// 变量节点97
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_97(
.clk(clk),
.rst(rst),
.initial_value(initial_value[97]),
.initial_value_enable(initial_value_enable[97]),
.initial_down(initial_down[97]),
.check_value_input(value_check_to_variable_97),
.check_enable_input(enable_check_to_variable_97),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_97_to_decision),
.value_variable_to_check(value_variable_97_to_check),
.variable_enable(enable_variable_97_to_check)
);

// 变量节点98
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_98(
.clk(clk),
.rst(rst),
.initial_value(initial_value[98]),
.initial_value_enable(initial_value_enable[98]),
.initial_down(initial_down[98]),
.check_value_input(value_check_to_variable_98),
.check_enable_input(enable_check_to_variable_98),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_98_to_decision),
.value_variable_to_check(value_variable_98_to_check),
.variable_enable(enable_variable_98_to_check)
);

// 变量节点99
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_99(
.clk(clk),
.rst(rst),
.initial_value(initial_value[99]),
.initial_value_enable(initial_value_enable[99]),
.initial_down(initial_down[99]),
.check_value_input(value_check_to_variable_99),
.check_enable_input(enable_check_to_variable_99),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_99_to_decision),
.value_variable_to_check(value_variable_99_to_check),
.variable_enable(enable_variable_99_to_check)
);

// 变量节点100
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_100(
.clk(clk),
.rst(rst),
.initial_value(initial_value[100]),
.initial_value_enable(initial_value_enable[100]),
.initial_down(initial_down[100]),
.check_value_input(value_check_to_variable_100),
.check_enable_input(enable_check_to_variable_100),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_100_to_decision),
.value_variable_to_check(value_variable_100_to_check),
.variable_enable(enable_variable_100_to_check)
);

// 变量节点101
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_101(
.clk(clk),
.rst(rst),
.initial_value(initial_value[101]),
.initial_value_enable(initial_value_enable[101]),
.initial_down(initial_down[101]),
.check_value_input(value_check_to_variable_101),
.check_enable_input(enable_check_to_variable_101),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_101_to_decision),
.value_variable_to_check(value_variable_101_to_check),
.variable_enable(enable_variable_101_to_check)
);

// 变量节点102
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_102(
.clk(clk),
.rst(rst),
.initial_value(initial_value[102]),
.initial_value_enable(initial_value_enable[102]),
.initial_down(initial_down[102]),
.check_value_input(value_check_to_variable_102),
.check_enable_input(enable_check_to_variable_102),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_102_to_decision),
.value_variable_to_check(value_variable_102_to_check),
.variable_enable(enable_variable_102_to_check)
);

// 变量节点103
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_103(
.clk(clk),
.rst(rst),
.initial_value(initial_value[103]),
.initial_value_enable(initial_value_enable[103]),
.initial_down(initial_down[103]),
.check_value_input(value_check_to_variable_103),
.check_enable_input(enable_check_to_variable_103),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_103_to_decision),
.value_variable_to_check(value_variable_103_to_check),
.variable_enable(enable_variable_103_to_check)
);

// 变量节点104
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_104(
.clk(clk),
.rst(rst),
.initial_value(initial_value[104]),
.initial_value_enable(initial_value_enable[104]),
.initial_down(initial_down[104]),
.check_value_input(value_check_to_variable_104),
.check_enable_input(enable_check_to_variable_104),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_104_to_decision),
.value_variable_to_check(value_variable_104_to_check),
.variable_enable(enable_variable_104_to_check)
);

// 变量节点105
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_105(
.clk(clk),
.rst(rst),
.initial_value(initial_value[105]),
.initial_value_enable(initial_value_enable[105]),
.initial_down(initial_down[105]),
.check_value_input(value_check_to_variable_105),
.check_enable_input(enable_check_to_variable_105),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_105_to_decision),
.value_variable_to_check(value_variable_105_to_check),
.variable_enable(enable_variable_105_to_check)
);

// 变量节点106
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_106(
.clk(clk),
.rst(rst),
.initial_value(initial_value[106]),
.initial_value_enable(initial_value_enable[106]),
.initial_down(initial_down[106]),
.check_value_input(value_check_to_variable_106),
.check_enable_input(enable_check_to_variable_106),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_106_to_decision),
.value_variable_to_check(value_variable_106_to_check),
.variable_enable(enable_variable_106_to_check)
);

// 变量节点107
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_107(
.clk(clk),
.rst(rst),
.initial_value(initial_value[107]),
.initial_value_enable(initial_value_enable[107]),
.initial_down(initial_down[107]),
.check_value_input(value_check_to_variable_107),
.check_enable_input(enable_check_to_variable_107),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_107_to_decision),
.value_variable_to_check(value_variable_107_to_check),
.variable_enable(enable_variable_107_to_check)
);

// 变量节点108
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_108(
.clk(clk),
.rst(rst),
.initial_value(initial_value[108]),
.initial_value_enable(initial_value_enable[108]),
.initial_down(initial_down[108]),
.check_value_input(value_check_to_variable_108),
.check_enable_input(enable_check_to_variable_108),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_108_to_decision),
.value_variable_to_check(value_variable_108_to_check),
.variable_enable(enable_variable_108_to_check)
);

// 变量节点109
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_109(
.clk(clk),
.rst(rst),
.initial_value(initial_value[109]),
.initial_value_enable(initial_value_enable[109]),
.initial_down(initial_down[109]),
.check_value_input(value_check_to_variable_109),
.check_enable_input(enable_check_to_variable_109),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_109_to_decision),
.value_variable_to_check(value_variable_109_to_check),
.variable_enable(enable_variable_109_to_check)
);

// 变量节点110
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_110(
.clk(clk),
.rst(rst),
.initial_value(initial_value[110]),
.initial_value_enable(initial_value_enable[110]),
.initial_down(initial_down[110]),
.check_value_input(value_check_to_variable_110),
.check_enable_input(enable_check_to_variable_110),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_110_to_decision),
.value_variable_to_check(value_variable_110_to_check),
.variable_enable(enable_variable_110_to_check)
);

// 变量节点111
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_111(
.clk(clk),
.rst(rst),
.initial_value(initial_value[111]),
.initial_value_enable(initial_value_enable[111]),
.initial_down(initial_down[111]),
.check_value_input(value_check_to_variable_111),
.check_enable_input(enable_check_to_variable_111),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_111_to_decision),
.value_variable_to_check(value_variable_111_to_check),
.variable_enable(enable_variable_111_to_check)
);

// 变量节点112
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_112(
.clk(clk),
.rst(rst),
.initial_value(initial_value[112]),
.initial_value_enable(initial_value_enable[112]),
.initial_down(initial_down[112]),
.check_value_input(value_check_to_variable_112),
.check_enable_input(enable_check_to_variable_112),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_112_to_decision),
.value_variable_to_check(value_variable_112_to_check),
.variable_enable(enable_variable_112_to_check)
);

// 变量节点113
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_113(
.clk(clk),
.rst(rst),
.initial_value(initial_value[113]),
.initial_value_enable(initial_value_enable[113]),
.initial_down(initial_down[113]),
.check_value_input(value_check_to_variable_113),
.check_enable_input(enable_check_to_variable_113),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_113_to_decision),
.value_variable_to_check(value_variable_113_to_check),
.variable_enable(enable_variable_113_to_check)
);

// 变量节点114
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_114(
.clk(clk),
.rst(rst),
.initial_value(initial_value[114]),
.initial_value_enable(initial_value_enable[114]),
.initial_down(initial_down[114]),
.check_value_input(value_check_to_variable_114),
.check_enable_input(enable_check_to_variable_114),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_114_to_decision),
.value_variable_to_check(value_variable_114_to_check),
.variable_enable(enable_variable_114_to_check)
);

// 变量节点115
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_115(
.clk(clk),
.rst(rst),
.initial_value(initial_value[115]),
.initial_value_enable(initial_value_enable[115]),
.initial_down(initial_down[115]),
.check_value_input(value_check_to_variable_115),
.check_enable_input(enable_check_to_variable_115),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_115_to_decision),
.value_variable_to_check(value_variable_115_to_check),
.variable_enable(enable_variable_115_to_check)
);

// 变量节点116
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_116(
.clk(clk),
.rst(rst),
.initial_value(initial_value[116]),
.initial_value_enable(initial_value_enable[116]),
.initial_down(initial_down[116]),
.check_value_input(value_check_to_variable_116),
.check_enable_input(enable_check_to_variable_116),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_116_to_decision),
.value_variable_to_check(value_variable_116_to_check),
.variable_enable(enable_variable_116_to_check)
);

// 变量节点117
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_117(
.clk(clk),
.rst(rst),
.initial_value(initial_value[117]),
.initial_value_enable(initial_value_enable[117]),
.initial_down(initial_down[117]),
.check_value_input(value_check_to_variable_117),
.check_enable_input(enable_check_to_variable_117),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_117_to_decision),
.value_variable_to_check(value_variable_117_to_check),
.variable_enable(enable_variable_117_to_check)
);

// 变量节点118
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_118(
.clk(clk),
.rst(rst),
.initial_value(initial_value[118]),
.initial_value_enable(initial_value_enable[118]),
.initial_down(initial_down[118]),
.check_value_input(value_check_to_variable_118),
.check_enable_input(enable_check_to_variable_118),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_118_to_decision),
.value_variable_to_check(value_variable_118_to_check),
.variable_enable(enable_variable_118_to_check)
);

// 变量节点119
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_119(
.clk(clk),
.rst(rst),
.initial_value(initial_value[119]),
.initial_value_enable(initial_value_enable[119]),
.initial_down(initial_down[119]),
.check_value_input(value_check_to_variable_119),
.check_enable_input(enable_check_to_variable_119),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_119_to_decision),
.value_variable_to_check(value_variable_119_to_check),
.variable_enable(enable_variable_119_to_check)
);

// 变量节点120
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_120(
.clk(clk),
.rst(rst),
.initial_value(initial_value[120]),
.initial_value_enable(initial_value_enable[120]),
.initial_down(initial_down[120]),
.check_value_input(value_check_to_variable_120),
.check_enable_input(enable_check_to_variable_120),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_120_to_decision),
.value_variable_to_check(value_variable_120_to_check),
.variable_enable(enable_variable_120_to_check)
);

// 变量节点121
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_121(
.clk(clk),
.rst(rst),
.initial_value(initial_value[121]),
.initial_value_enable(initial_value_enable[121]),
.initial_down(initial_down[121]),
.check_value_input(value_check_to_variable_121),
.check_enable_input(enable_check_to_variable_121),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_121_to_decision),
.value_variable_to_check(value_variable_121_to_check),
.variable_enable(enable_variable_121_to_check)
);

// 变量节点122
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_122(
.clk(clk),
.rst(rst),
.initial_value(initial_value[122]),
.initial_value_enable(initial_value_enable[122]),
.initial_down(initial_down[122]),
.check_value_input(value_check_to_variable_122),
.check_enable_input(enable_check_to_variable_122),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_122_to_decision),
.value_variable_to_check(value_variable_122_to_check),
.variable_enable(enable_variable_122_to_check)
);

// 变量节点123
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_123(
.clk(clk),
.rst(rst),
.initial_value(initial_value[123]),
.initial_value_enable(initial_value_enable[123]),
.initial_down(initial_down[123]),
.check_value_input(value_check_to_variable_123),
.check_enable_input(enable_check_to_variable_123),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_123_to_decision),
.value_variable_to_check(value_variable_123_to_check),
.variable_enable(enable_variable_123_to_check)
);

// 变量节点124
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_124(
.clk(clk),
.rst(rst),
.initial_value(initial_value[124]),
.initial_value_enable(initial_value_enable[124]),
.initial_down(initial_down[124]),
.check_value_input(value_check_to_variable_124),
.check_enable_input(enable_check_to_variable_124),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_124_to_decision),
.value_variable_to_check(value_variable_124_to_check),
.variable_enable(enable_variable_124_to_check)
);

// 变量节点125
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_125(
.clk(clk),
.rst(rst),
.initial_value(initial_value[125]),
.initial_value_enable(initial_value_enable[125]),
.initial_down(initial_down[125]),
.check_value_input(value_check_to_variable_125),
.check_enable_input(enable_check_to_variable_125),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_125_to_decision),
.value_variable_to_check(value_variable_125_to_check),
.variable_enable(enable_variable_125_to_check)
);

// 变量节点126
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_126(
.clk(clk),
.rst(rst),
.initial_value(initial_value[126]),
.initial_value_enable(initial_value_enable[126]),
.initial_down(initial_down[126]),
.check_value_input(value_check_to_variable_126),
.check_enable_input(enable_check_to_variable_126),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_126_to_decision),
.value_variable_to_check(value_variable_126_to_check),
.variable_enable(enable_variable_126_to_check)
);

// 变量节点127
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_127(
.clk(clk),
.rst(rst),
.initial_value(initial_value[127]),
.initial_value_enable(initial_value_enable[127]),
.initial_down(initial_down[127]),
.check_value_input(value_check_to_variable_127),
.check_enable_input(enable_check_to_variable_127),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_127_to_decision),
.value_variable_to_check(value_variable_127_to_check),
.variable_enable(enable_variable_127_to_check)
);

// 变量节点128
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_128(
.clk(clk),
.rst(rst),
.initial_value(initial_value[128]),
.initial_value_enable(initial_value_enable[128]),
.initial_down(initial_down[128]),
.check_value_input(value_check_to_variable_128),
.check_enable_input(enable_check_to_variable_128),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_128_to_decision),
.value_variable_to_check(value_variable_128_to_check),
.variable_enable(enable_variable_128_to_check)
);

// 变量节点129
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_129(
.clk(clk),
.rst(rst),
.initial_value(initial_value[129]),
.initial_value_enable(initial_value_enable[129]),
.initial_down(initial_down[129]),
.check_value_input(value_check_to_variable_129),
.check_enable_input(enable_check_to_variable_129),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_129_to_decision),
.value_variable_to_check(value_variable_129_to_check),
.variable_enable(enable_variable_129_to_check)
);

// 变量节点130
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_130(
.clk(clk),
.rst(rst),
.initial_value(initial_value[130]),
.initial_value_enable(initial_value_enable[130]),
.initial_down(initial_down[130]),
.check_value_input(value_check_to_variable_130),
.check_enable_input(enable_check_to_variable_130),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_130_to_decision),
.value_variable_to_check(value_variable_130_to_check),
.variable_enable(enable_variable_130_to_check)
);

// 变量节点131
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_131(
.clk(clk),
.rst(rst),
.initial_value(initial_value[131]),
.initial_value_enable(initial_value_enable[131]),
.initial_down(initial_down[131]),
.check_value_input(value_check_to_variable_131),
.check_enable_input(enable_check_to_variable_131),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_131_to_decision),
.value_variable_to_check(value_variable_131_to_check),
.variable_enable(enable_variable_131_to_check)
);

// 变量节点132
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_132(
.clk(clk),
.rst(rst),
.initial_value(initial_value[132]),
.initial_value_enable(initial_value_enable[132]),
.initial_down(initial_down[132]),
.check_value_input(value_check_to_variable_132),
.check_enable_input(enable_check_to_variable_132),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_132_to_decision),
.value_variable_to_check(value_variable_132_to_check),
.variable_enable(enable_variable_132_to_check)
);

// 变量节点133
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_133(
.clk(clk),
.rst(rst),
.initial_value(initial_value[133]),
.initial_value_enable(initial_value_enable[133]),
.initial_down(initial_down[133]),
.check_value_input(value_check_to_variable_133),
.check_enable_input(enable_check_to_variable_133),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_133_to_decision),
.value_variable_to_check(value_variable_133_to_check),
.variable_enable(enable_variable_133_to_check)
);

// 变量节点134
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_134(
.clk(clk),
.rst(rst),
.initial_value(initial_value[134]),
.initial_value_enable(initial_value_enable[134]),
.initial_down(initial_down[134]),
.check_value_input(value_check_to_variable_134),
.check_enable_input(enable_check_to_variable_134),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_134_to_decision),
.value_variable_to_check(value_variable_134_to_check),
.variable_enable(enable_variable_134_to_check)
);

// 变量节点135
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_135(
.clk(clk),
.rst(rst),
.initial_value(initial_value[135]),
.initial_value_enable(initial_value_enable[135]),
.initial_down(initial_down[135]),
.check_value_input(value_check_to_variable_135),
.check_enable_input(enable_check_to_variable_135),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_135_to_decision),
.value_variable_to_check(value_variable_135_to_check),
.variable_enable(enable_variable_135_to_check)
);

// 变量节点136
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_136(
.clk(clk),
.rst(rst),
.initial_value(initial_value[136]),
.initial_value_enable(initial_value_enable[136]),
.initial_down(initial_down[136]),
.check_value_input(value_check_to_variable_136),
.check_enable_input(enable_check_to_variable_136),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_136_to_decision),
.value_variable_to_check(value_variable_136_to_check),
.variable_enable(enable_variable_136_to_check)
);

// 变量节点137
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_137(
.clk(clk),
.rst(rst),
.initial_value(initial_value[137]),
.initial_value_enable(initial_value_enable[137]),
.initial_down(initial_down[137]),
.check_value_input(value_check_to_variable_137),
.check_enable_input(enable_check_to_variable_137),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_137_to_decision),
.value_variable_to_check(value_variable_137_to_check),
.variable_enable(enable_variable_137_to_check)
);

// 变量节点138
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_138(
.clk(clk),
.rst(rst),
.initial_value(initial_value[138]),
.initial_value_enable(initial_value_enable[138]),
.initial_down(initial_down[138]),
.check_value_input(value_check_to_variable_138),
.check_enable_input(enable_check_to_variable_138),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_138_to_decision),
.value_variable_to_check(value_variable_138_to_check),
.variable_enable(enable_variable_138_to_check)
);

// 变量节点139
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_139(
.clk(clk),
.rst(rst),
.initial_value(initial_value[139]),
.initial_value_enable(initial_value_enable[139]),
.initial_down(initial_down[139]),
.check_value_input(value_check_to_variable_139),
.check_enable_input(enable_check_to_variable_139),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_139_to_decision),
.value_variable_to_check(value_variable_139_to_check),
.variable_enable(enable_variable_139_to_check)
);

// 变量节点140
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_140(
.clk(clk),
.rst(rst),
.initial_value(initial_value[140]),
.initial_value_enable(initial_value_enable[140]),
.initial_down(initial_down[140]),
.check_value_input(value_check_to_variable_140),
.check_enable_input(enable_check_to_variable_140),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_140_to_decision),
.value_variable_to_check(value_variable_140_to_check),
.variable_enable(enable_variable_140_to_check)
);

// 变量节点141
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_141(
.clk(clk),
.rst(rst),
.initial_value(initial_value[141]),
.initial_value_enable(initial_value_enable[141]),
.initial_down(initial_down[141]),
.check_value_input(value_check_to_variable_141),
.check_enable_input(enable_check_to_variable_141),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_141_to_decision),
.value_variable_to_check(value_variable_141_to_check),
.variable_enable(enable_variable_141_to_check)
);

// 变量节点142
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_142(
.clk(clk),
.rst(rst),
.initial_value(initial_value[142]),
.initial_value_enable(initial_value_enable[142]),
.initial_down(initial_down[142]),
.check_value_input(value_check_to_variable_142),
.check_enable_input(enable_check_to_variable_142),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_142_to_decision),
.value_variable_to_check(value_variable_142_to_check),
.variable_enable(enable_variable_142_to_check)
);

// 变量节点143
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_143(
.clk(clk),
.rst(rst),
.initial_value(initial_value[143]),
.initial_value_enable(initial_value_enable[143]),
.initial_down(initial_down[143]),
.check_value_input(value_check_to_variable_143),
.check_enable_input(enable_check_to_variable_143),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_143_to_decision),
.value_variable_to_check(value_variable_143_to_check),
.variable_enable(enable_variable_143_to_check)
);

// 变量节点144
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_144(
.clk(clk),
.rst(rst),
.initial_value(initial_value[144]),
.initial_value_enable(initial_value_enable[144]),
.initial_down(initial_down[144]),
.check_value_input(value_check_to_variable_144),
.check_enable_input(enable_check_to_variable_144),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_144_to_decision),
.value_variable_to_check(value_variable_144_to_check),
.variable_enable(enable_variable_144_to_check)
);

// 变量节点145
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_145(
.clk(clk),
.rst(rst),
.initial_value(initial_value[145]),
.initial_value_enable(initial_value_enable[145]),
.initial_down(initial_down[145]),
.check_value_input(value_check_to_variable_145),
.check_enable_input(enable_check_to_variable_145),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_145_to_decision),
.value_variable_to_check(value_variable_145_to_check),
.variable_enable(enable_variable_145_to_check)
);

// 变量节点146
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_146(
.clk(clk),
.rst(rst),
.initial_value(initial_value[146]),
.initial_value_enable(initial_value_enable[146]),
.initial_down(initial_down[146]),
.check_value_input(value_check_to_variable_146),
.check_enable_input(enable_check_to_variable_146),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_146_to_decision),
.value_variable_to_check(value_variable_146_to_check),
.variable_enable(enable_variable_146_to_check)
);

// 变量节点147
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_147(
.clk(clk),
.rst(rst),
.initial_value(initial_value[147]),
.initial_value_enable(initial_value_enable[147]),
.initial_down(initial_down[147]),
.check_value_input(value_check_to_variable_147),
.check_enable_input(enable_check_to_variable_147),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_147_to_decision),
.value_variable_to_check(value_variable_147_to_check),
.variable_enable(enable_variable_147_to_check)
);

// 变量节点148
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_148(
.clk(clk),
.rst(rst),
.initial_value(initial_value[148]),
.initial_value_enable(initial_value_enable[148]),
.initial_down(initial_down[148]),
.check_value_input(value_check_to_variable_148),
.check_enable_input(enable_check_to_variable_148),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_148_to_decision),
.value_variable_to_check(value_variable_148_to_check),
.variable_enable(enable_variable_148_to_check)
);

// 变量节点149
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_149(
.clk(clk),
.rst(rst),
.initial_value(initial_value[149]),
.initial_value_enable(initial_value_enable[149]),
.initial_down(initial_down[149]),
.check_value_input(value_check_to_variable_149),
.check_enable_input(enable_check_to_variable_149),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_149_to_decision),
.value_variable_to_check(value_variable_149_to_check),
.variable_enable(enable_variable_149_to_check)
);

// 变量节点150
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_150(
.clk(clk),
.rst(rst),
.initial_value(initial_value[150]),
.initial_value_enable(initial_value_enable[150]),
.initial_down(initial_down[150]),
.check_value_input(value_check_to_variable_150),
.check_enable_input(enable_check_to_variable_150),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_150_to_decision),
.value_variable_to_check(value_variable_150_to_check),
.variable_enable(enable_variable_150_to_check)
);

// 变量节点151
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_151(
.clk(clk),
.rst(rst),
.initial_value(initial_value[151]),
.initial_value_enable(initial_value_enable[151]),
.initial_down(initial_down[151]),
.check_value_input(value_check_to_variable_151),
.check_enable_input(enable_check_to_variable_151),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_151_to_decision),
.value_variable_to_check(value_variable_151_to_check),
.variable_enable(enable_variable_151_to_check)
);

// 变量节点152
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_152(
.clk(clk),
.rst(rst),
.initial_value(initial_value[152]),
.initial_value_enable(initial_value_enable[152]),
.initial_down(initial_down[152]),
.check_value_input(value_check_to_variable_152),
.check_enable_input(enable_check_to_variable_152),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_152_to_decision),
.value_variable_to_check(value_variable_152_to_check),
.variable_enable(enable_variable_152_to_check)
);

// 变量节点153
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_153(
.clk(clk),
.rst(rst),
.initial_value(initial_value[153]),
.initial_value_enable(initial_value_enable[153]),
.initial_down(initial_down[153]),
.check_value_input(value_check_to_variable_153),
.check_enable_input(enable_check_to_variable_153),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_153_to_decision),
.value_variable_to_check(value_variable_153_to_check),
.variable_enable(enable_variable_153_to_check)
);

// 变量节点154
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_154(
.clk(clk),
.rst(rst),
.initial_value(initial_value[154]),
.initial_value_enable(initial_value_enable[154]),
.initial_down(initial_down[154]),
.check_value_input(value_check_to_variable_154),
.check_enable_input(enable_check_to_variable_154),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_154_to_decision),
.value_variable_to_check(value_variable_154_to_check),
.variable_enable(enable_variable_154_to_check)
);

// 变量节点155
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_155(
.clk(clk),
.rst(rst),
.initial_value(initial_value[155]),
.initial_value_enable(initial_value_enable[155]),
.initial_down(initial_down[155]),
.check_value_input(value_check_to_variable_155),
.check_enable_input(enable_check_to_variable_155),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_155_to_decision),
.value_variable_to_check(value_variable_155_to_check),
.variable_enable(enable_variable_155_to_check)
);

// 变量节点156
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_156(
.clk(clk),
.rst(rst),
.initial_value(initial_value[156]),
.initial_value_enable(initial_value_enable[156]),
.initial_down(initial_down[156]),
.check_value_input(value_check_to_variable_156),
.check_enable_input(enable_check_to_variable_156),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_156_to_decision),
.value_variable_to_check(value_variable_156_to_check),
.variable_enable(enable_variable_156_to_check)
);

// 变量节点157
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_157(
.clk(clk),
.rst(rst),
.initial_value(initial_value[157]),
.initial_value_enable(initial_value_enable[157]),
.initial_down(initial_down[157]),
.check_value_input(value_check_to_variable_157),
.check_enable_input(enable_check_to_variable_157),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_157_to_decision),
.value_variable_to_check(value_variable_157_to_check),
.variable_enable(enable_variable_157_to_check)
);

// 变量节点158
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_158(
.clk(clk),
.rst(rst),
.initial_value(initial_value[158]),
.initial_value_enable(initial_value_enable[158]),
.initial_down(initial_down[158]),
.check_value_input(value_check_to_variable_158),
.check_enable_input(enable_check_to_variable_158),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_158_to_decision),
.value_variable_to_check(value_variable_158_to_check),
.variable_enable(enable_variable_158_to_check)
);

// 变量节点159
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_159(
.clk(clk),
.rst(rst),
.initial_value(initial_value[159]),
.initial_value_enable(initial_value_enable[159]),
.initial_down(initial_down[159]),
.check_value_input(value_check_to_variable_159),
.check_enable_input(enable_check_to_variable_159),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_159_to_decision),
.value_variable_to_check(value_variable_159_to_check),
.variable_enable(enable_variable_159_to_check)
);

// 变量节点160
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_160(
.clk(clk),
.rst(rst),
.initial_value(initial_value[160]),
.initial_value_enable(initial_value_enable[160]),
.initial_down(initial_down[160]),
.check_value_input(value_check_to_variable_160),
.check_enable_input(enable_check_to_variable_160),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_160_to_decision),
.value_variable_to_check(value_variable_160_to_check),
.variable_enable(enable_variable_160_to_check)
);

// 变量节点161
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_161(
.clk(clk),
.rst(rst),
.initial_value(initial_value[161]),
.initial_value_enable(initial_value_enable[161]),
.initial_down(initial_down[161]),
.check_value_input(value_check_to_variable_161),
.check_enable_input(enable_check_to_variable_161),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_161_to_decision),
.value_variable_to_check(value_variable_161_to_check),
.variable_enable(enable_variable_161_to_check)
);

// 变量节点162
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_162(
.clk(clk),
.rst(rst),
.initial_value(initial_value[162]),
.initial_value_enable(initial_value_enable[162]),
.initial_down(initial_down[162]),
.check_value_input(value_check_to_variable_162),
.check_enable_input(enable_check_to_variable_162),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_162_to_decision),
.value_variable_to_check(value_variable_162_to_check),
.variable_enable(enable_variable_162_to_check)
);

// 变量节点163
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_163(
.clk(clk),
.rst(rst),
.initial_value(initial_value[163]),
.initial_value_enable(initial_value_enable[163]),
.initial_down(initial_down[163]),
.check_value_input(value_check_to_variable_163),
.check_enable_input(enable_check_to_variable_163),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_163_to_decision),
.value_variable_to_check(value_variable_163_to_check),
.variable_enable(enable_variable_163_to_check)
);

// 变量节点164
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_164(
.clk(clk),
.rst(rst),
.initial_value(initial_value[164]),
.initial_value_enable(initial_value_enable[164]),
.initial_down(initial_down[164]),
.check_value_input(value_check_to_variable_164),
.check_enable_input(enable_check_to_variable_164),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_164_to_decision),
.value_variable_to_check(value_variable_164_to_check),
.variable_enable(enable_variable_164_to_check)
);

// 变量节点165
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_165(
.clk(clk),
.rst(rst),
.initial_value(initial_value[165]),
.initial_value_enable(initial_value_enable[165]),
.initial_down(initial_down[165]),
.check_value_input(value_check_to_variable_165),
.check_enable_input(enable_check_to_variable_165),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_165_to_decision),
.value_variable_to_check(value_variable_165_to_check),
.variable_enable(enable_variable_165_to_check)
);

// 变量节点166
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_166(
.clk(clk),
.rst(rst),
.initial_value(initial_value[166]),
.initial_value_enable(initial_value_enable[166]),
.initial_down(initial_down[166]),
.check_value_input(value_check_to_variable_166),
.check_enable_input(enable_check_to_variable_166),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_166_to_decision),
.value_variable_to_check(value_variable_166_to_check),
.variable_enable(enable_variable_166_to_check)
);

// 变量节点167
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_167(
.clk(clk),
.rst(rst),
.initial_value(initial_value[167]),
.initial_value_enable(initial_value_enable[167]),
.initial_down(initial_down[167]),
.check_value_input(value_check_to_variable_167),
.check_enable_input(enable_check_to_variable_167),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_167_to_decision),
.value_variable_to_check(value_variable_167_to_check),
.variable_enable(enable_variable_167_to_check)
);

// 变量节点168
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_168(
.clk(clk),
.rst(rst),
.initial_value(initial_value[168]),
.initial_value_enable(initial_value_enable[168]),
.initial_down(initial_down[168]),
.check_value_input(value_check_to_variable_168),
.check_enable_input(enable_check_to_variable_168),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_168_to_decision),
.value_variable_to_check(value_variable_168_to_check),
.variable_enable(enable_variable_168_to_check)
);

// 变量节点169
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_169(
.clk(clk),
.rst(rst),
.initial_value(initial_value[169]),
.initial_value_enable(initial_value_enable[169]),
.initial_down(initial_down[169]),
.check_value_input(value_check_to_variable_169),
.check_enable_input(enable_check_to_variable_169),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_169_to_decision),
.value_variable_to_check(value_variable_169_to_check),
.variable_enable(enable_variable_169_to_check)
);

// 变量节点170
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_170(
.clk(clk),
.rst(rst),
.initial_value(initial_value[170]),
.initial_value_enable(initial_value_enable[170]),
.initial_down(initial_down[170]),
.check_value_input(value_check_to_variable_170),
.check_enable_input(enable_check_to_variable_170),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_170_to_decision),
.value_variable_to_check(value_variable_170_to_check),
.variable_enable(enable_variable_170_to_check)
);

// 变量节点171
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_171(
.clk(clk),
.rst(rst),
.initial_value(initial_value[171]),
.initial_value_enable(initial_value_enable[171]),
.initial_down(initial_down[171]),
.check_value_input(value_check_to_variable_171),
.check_enable_input(enable_check_to_variable_171),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_171_to_decision),
.value_variable_to_check(value_variable_171_to_check),
.variable_enable(enable_variable_171_to_check)
);

// 变量节点172
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_172(
.clk(clk),
.rst(rst),
.initial_value(initial_value[172]),
.initial_value_enable(initial_value_enable[172]),
.initial_down(initial_down[172]),
.check_value_input(value_check_to_variable_172),
.check_enable_input(enable_check_to_variable_172),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_172_to_decision),
.value_variable_to_check(value_variable_172_to_check),
.variable_enable(enable_variable_172_to_check)
);

// 变量节点173
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_173(
.clk(clk),
.rst(rst),
.initial_value(initial_value[173]),
.initial_value_enable(initial_value_enable[173]),
.initial_down(initial_down[173]),
.check_value_input(value_check_to_variable_173),
.check_enable_input(enable_check_to_variable_173),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_173_to_decision),
.value_variable_to_check(value_variable_173_to_check),
.variable_enable(enable_variable_173_to_check)
);

// 变量节点174
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_174(
.clk(clk),
.rst(rst),
.initial_value(initial_value[174]),
.initial_value_enable(initial_value_enable[174]),
.initial_down(initial_down[174]),
.check_value_input(value_check_to_variable_174),
.check_enable_input(enable_check_to_variable_174),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_174_to_decision),
.value_variable_to_check(value_variable_174_to_check),
.variable_enable(enable_variable_174_to_check)
);

// 变量节点175
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_175(
.clk(clk),
.rst(rst),
.initial_value(initial_value[175]),
.initial_value_enable(initial_value_enable[175]),
.initial_down(initial_down[175]),
.check_value_input(value_check_to_variable_175),
.check_enable_input(enable_check_to_variable_175),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_175_to_decision),
.value_variable_to_check(value_variable_175_to_check),
.variable_enable(enable_variable_175_to_check)
);

// 变量节点176
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_176(
.clk(clk),
.rst(rst),
.initial_value(initial_value[176]),
.initial_value_enable(initial_value_enable[176]),
.initial_down(initial_down[176]),
.check_value_input(value_check_to_variable_176),
.check_enable_input(enable_check_to_variable_176),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_176_to_decision),
.value_variable_to_check(value_variable_176_to_check),
.variable_enable(enable_variable_176_to_check)
);

// 变量节点177
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_177(
.clk(clk),
.rst(rst),
.initial_value(initial_value[177]),
.initial_value_enable(initial_value_enable[177]),
.initial_down(initial_down[177]),
.check_value_input(value_check_to_variable_177),
.check_enable_input(enable_check_to_variable_177),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_177_to_decision),
.value_variable_to_check(value_variable_177_to_check),
.variable_enable(enable_variable_177_to_check)
);

// 变量节点178
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_178(
.clk(clk),
.rst(rst),
.initial_value(initial_value[178]),
.initial_value_enable(initial_value_enable[178]),
.initial_down(initial_down[178]),
.check_value_input(value_check_to_variable_178),
.check_enable_input(enable_check_to_variable_178),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_178_to_decision),
.value_variable_to_check(value_variable_178_to_check),
.variable_enable(enable_variable_178_to_check)
);

// 变量节点179
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_179(
.clk(clk),
.rst(rst),
.initial_value(initial_value[179]),
.initial_value_enable(initial_value_enable[179]),
.initial_down(initial_down[179]),
.check_value_input(value_check_to_variable_179),
.check_enable_input(enable_check_to_variable_179),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_179_to_decision),
.value_variable_to_check(value_variable_179_to_check),
.variable_enable(enable_variable_179_to_check)
);

// 变量节点180
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_180(
.clk(clk),
.rst(rst),
.initial_value(initial_value[180]),
.initial_value_enable(initial_value_enable[180]),
.initial_down(initial_down[180]),
.check_value_input(value_check_to_variable_180),
.check_enable_input(enable_check_to_variable_180),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_180_to_decision),
.value_variable_to_check(value_variable_180_to_check),
.variable_enable(enable_variable_180_to_check)
);

// 变量节点181
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_181(
.clk(clk),
.rst(rst),
.initial_value(initial_value[181]),
.initial_value_enable(initial_value_enable[181]),
.initial_down(initial_down[181]),
.check_value_input(value_check_to_variable_181),
.check_enable_input(enable_check_to_variable_181),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_181_to_decision),
.value_variable_to_check(value_variable_181_to_check),
.variable_enable(enable_variable_181_to_check)
);

// 变量节点182
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_182(
.clk(clk),
.rst(rst),
.initial_value(initial_value[182]),
.initial_value_enable(initial_value_enable[182]),
.initial_down(initial_down[182]),
.check_value_input(value_check_to_variable_182),
.check_enable_input(enable_check_to_variable_182),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_182_to_decision),
.value_variable_to_check(value_variable_182_to_check),
.variable_enable(enable_variable_182_to_check)
);

// 变量节点183
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_183(
.clk(clk),
.rst(rst),
.initial_value(initial_value[183]),
.initial_value_enable(initial_value_enable[183]),
.initial_down(initial_down[183]),
.check_value_input(value_check_to_variable_183),
.check_enable_input(enable_check_to_variable_183),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_183_to_decision),
.value_variable_to_check(value_variable_183_to_check),
.variable_enable(enable_variable_183_to_check)
);

// 变量节点184
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_184(
.clk(clk),
.rst(rst),
.initial_value(initial_value[184]),
.initial_value_enable(initial_value_enable[184]),
.initial_down(initial_down[184]),
.check_value_input(value_check_to_variable_184),
.check_enable_input(enable_check_to_variable_184),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_184_to_decision),
.value_variable_to_check(value_variable_184_to_check),
.variable_enable(enable_variable_184_to_check)
);

// 变量节点185
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_185(
.clk(clk),
.rst(rst),
.initial_value(initial_value[185]),
.initial_value_enable(initial_value_enable[185]),
.initial_down(initial_down[185]),
.check_value_input(value_check_to_variable_185),
.check_enable_input(enable_check_to_variable_185),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_185_to_decision),
.value_variable_to_check(value_variable_185_to_check),
.variable_enable(enable_variable_185_to_check)
);

// 变量节点186
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_186(
.clk(clk),
.rst(rst),
.initial_value(initial_value[186]),
.initial_value_enable(initial_value_enable[186]),
.initial_down(initial_down[186]),
.check_value_input(value_check_to_variable_186),
.check_enable_input(enable_check_to_variable_186),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_186_to_decision),
.value_variable_to_check(value_variable_186_to_check),
.variable_enable(enable_variable_186_to_check)
);

// 变量节点187
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_187(
.clk(clk),
.rst(rst),
.initial_value(initial_value[187]),
.initial_value_enable(initial_value_enable[187]),
.initial_down(initial_down[187]),
.check_value_input(value_check_to_variable_187),
.check_enable_input(enable_check_to_variable_187),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_187_to_decision),
.value_variable_to_check(value_variable_187_to_check),
.variable_enable(enable_variable_187_to_check)
);

// 变量节点188
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_188(
.clk(clk),
.rst(rst),
.initial_value(initial_value[188]),
.initial_value_enable(initial_value_enable[188]),
.initial_down(initial_down[188]),
.check_value_input(value_check_to_variable_188),
.check_enable_input(enable_check_to_variable_188),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_188_to_decision),
.value_variable_to_check(value_variable_188_to_check),
.variable_enable(enable_variable_188_to_check)
);

// 变量节点189
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_189(
.clk(clk),
.rst(rst),
.initial_value(initial_value[189]),
.initial_value_enable(initial_value_enable[189]),
.initial_down(initial_down[189]),
.check_value_input(value_check_to_variable_189),
.check_enable_input(enable_check_to_variable_189),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_189_to_decision),
.value_variable_to_check(value_variable_189_to_check),
.variable_enable(enable_variable_189_to_check)
);

// 变量节点190
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_190(
.clk(clk),
.rst(rst),
.initial_value(initial_value[190]),
.initial_value_enable(initial_value_enable[190]),
.initial_down(initial_down[190]),
.check_value_input(value_check_to_variable_190),
.check_enable_input(enable_check_to_variable_190),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_190_to_decision),
.value_variable_to_check(value_variable_190_to_check),
.variable_enable(enable_variable_190_to_check)
);

// 变量节点191
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_191(
.clk(clk),
.rst(rst),
.initial_value(initial_value[191]),
.initial_value_enable(initial_value_enable[191]),
.initial_down(initial_down[191]),
.check_value_input(value_check_to_variable_191),
.check_enable_input(enable_check_to_variable_191),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_191_to_decision),
.value_variable_to_check(value_variable_191_to_check),
.variable_enable(enable_variable_191_to_check)
);

// 变量节点192
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_192(
.clk(clk),
.rst(rst),
.initial_value(initial_value[192]),
.initial_value_enable(initial_value_enable[192]),
.initial_down(initial_down[192]),
.check_value_input(value_check_to_variable_192),
.check_enable_input(enable_check_to_variable_192),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_192_to_decision),
.value_variable_to_check(value_variable_192_to_check),
.variable_enable(enable_variable_192_to_check)
);

// 变量节点193
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_193(
.clk(clk),
.rst(rst),
.initial_value(initial_value[193]),
.initial_value_enable(initial_value_enable[193]),
.initial_down(initial_down[193]),
.check_value_input(value_check_to_variable_193),
.check_enable_input(enable_check_to_variable_193),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_193_to_decision),
.value_variable_to_check(value_variable_193_to_check),
.variable_enable(enable_variable_193_to_check)
);

// 变量节点194
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_194(
.clk(clk),
.rst(rst),
.initial_value(initial_value[194]),
.initial_value_enable(initial_value_enable[194]),
.initial_down(initial_down[194]),
.check_value_input(value_check_to_variable_194),
.check_enable_input(enable_check_to_variable_194),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_194_to_decision),
.value_variable_to_check(value_variable_194_to_check),
.variable_enable(enable_variable_194_to_check)
);

// 变量节点195
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_195(
.clk(clk),
.rst(rst),
.initial_value(initial_value[195]),
.initial_value_enable(initial_value_enable[195]),
.initial_down(initial_down[195]),
.check_value_input(value_check_to_variable_195),
.check_enable_input(enable_check_to_variable_195),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_195_to_decision),
.value_variable_to_check(value_variable_195_to_check),
.variable_enable(enable_variable_195_to_check)
);

// 变量节点196
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_196(
.clk(clk),
.rst(rst),
.initial_value(initial_value[196]),
.initial_value_enable(initial_value_enable[196]),
.initial_down(initial_down[196]),
.check_value_input(value_check_to_variable_196),
.check_enable_input(enable_check_to_variable_196),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_196_to_decision),
.value_variable_to_check(value_variable_196_to_check),
.variable_enable(enable_variable_196_to_check)
);

// 变量节点197
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_197(
.clk(clk),
.rst(rst),
.initial_value(initial_value[197]),
.initial_value_enable(initial_value_enable[197]),
.initial_down(initial_down[197]),
.check_value_input(value_check_to_variable_197),
.check_enable_input(enable_check_to_variable_197),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_197_to_decision),
.value_variable_to_check(value_variable_197_to_check),
.variable_enable(enable_variable_197_to_check)
);

// 变量节点198
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_198(
.clk(clk),
.rst(rst),
.initial_value(initial_value[198]),
.initial_value_enable(initial_value_enable[198]),
.initial_down(initial_down[198]),
.check_value_input(value_check_to_variable_198),
.check_enable_input(enable_check_to_variable_198),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_198_to_decision),
.value_variable_to_check(value_variable_198_to_check),
.variable_enable(enable_variable_198_to_check)
);

// 变量节点199
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_199(
.clk(clk),
.rst(rst),
.initial_value(initial_value[199]),
.initial_value_enable(initial_value_enable[199]),
.initial_down(initial_down[199]),
.check_value_input(value_check_to_variable_199),
.check_enable_input(enable_check_to_variable_199),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_199_to_decision),
.value_variable_to_check(value_variable_199_to_check),
.variable_enable(enable_variable_199_to_check)
);

// 变量节点200
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_200(
.clk(clk),
.rst(rst),
.initial_value(initial_value[200]),
.initial_value_enable(initial_value_enable[200]),
.initial_down(initial_down[200]),
.check_value_input(value_check_to_variable_200),
.check_enable_input(enable_check_to_variable_200),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_200_to_decision),
.value_variable_to_check(value_variable_200_to_check),
.variable_enable(enable_variable_200_to_check)
);

// 变量节点201
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_201(
.clk(clk),
.rst(rst),
.initial_value(initial_value[201]),
.initial_value_enable(initial_value_enable[201]),
.initial_down(initial_down[201]),
.check_value_input(value_check_to_variable_201),
.check_enable_input(enable_check_to_variable_201),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_201_to_decision),
.value_variable_to_check(value_variable_201_to_check),
.variable_enable(enable_variable_201_to_check)
);

// 变量节点202
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_202(
.clk(clk),
.rst(rst),
.initial_value(initial_value[202]),
.initial_value_enable(initial_value_enable[202]),
.initial_down(initial_down[202]),
.check_value_input(value_check_to_variable_202),
.check_enable_input(enable_check_to_variable_202),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_202_to_decision),
.value_variable_to_check(value_variable_202_to_check),
.variable_enable(enable_variable_202_to_check)
);

// 变量节点203
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_203(
.clk(clk),
.rst(rst),
.initial_value(initial_value[203]),
.initial_value_enable(initial_value_enable[203]),
.initial_down(initial_down[203]),
.check_value_input(value_check_to_variable_203),
.check_enable_input(enable_check_to_variable_203),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_203_to_decision),
.value_variable_to_check(value_variable_203_to_check),
.variable_enable(enable_variable_203_to_check)
);

// 变量节点204
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_204(
.clk(clk),
.rst(rst),
.initial_value(initial_value[204]),
.initial_value_enable(initial_value_enable[204]),
.initial_down(initial_down[204]),
.check_value_input(value_check_to_variable_204),
.check_enable_input(enable_check_to_variable_204),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_204_to_decision),
.value_variable_to_check(value_variable_204_to_check),
.variable_enable(enable_variable_204_to_check)
);

// 变量节点205
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_205(
.clk(clk),
.rst(rst),
.initial_value(initial_value[205]),
.initial_value_enable(initial_value_enable[205]),
.initial_down(initial_down[205]),
.check_value_input(value_check_to_variable_205),
.check_enable_input(enable_check_to_variable_205),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_205_to_decision),
.value_variable_to_check(value_variable_205_to_check),
.variable_enable(enable_variable_205_to_check)
);

// 变量节点206
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_206(
.clk(clk),
.rst(rst),
.initial_value(initial_value[206]),
.initial_value_enable(initial_value_enable[206]),
.initial_down(initial_down[206]),
.check_value_input(value_check_to_variable_206),
.check_enable_input(enable_check_to_variable_206),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_206_to_decision),
.value_variable_to_check(value_variable_206_to_check),
.variable_enable(enable_variable_206_to_check)
);

// 变量节点207
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_207(
.clk(clk),
.rst(rst),
.initial_value(initial_value[207]),
.initial_value_enable(initial_value_enable[207]),
.initial_down(initial_down[207]),
.check_value_input(value_check_to_variable_207),
.check_enable_input(enable_check_to_variable_207),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_207_to_decision),
.value_variable_to_check(value_variable_207_to_check),
.variable_enable(enable_variable_207_to_check)
);

// 变量节点208
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_208(
.clk(clk),
.rst(rst),
.initial_value(initial_value[208]),
.initial_value_enable(initial_value_enable[208]),
.initial_down(initial_down[208]),
.check_value_input(value_check_to_variable_208),
.check_enable_input(enable_check_to_variable_208),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_208_to_decision),
.value_variable_to_check(value_variable_208_to_check),
.variable_enable(enable_variable_208_to_check)
);

// 变量节点209
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_209(
.clk(clk),
.rst(rst),
.initial_value(initial_value[209]),
.initial_value_enable(initial_value_enable[209]),
.initial_down(initial_down[209]),
.check_value_input(value_check_to_variable_209),
.check_enable_input(enable_check_to_variable_209),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_209_to_decision),
.value_variable_to_check(value_variable_209_to_check),
.variable_enable(enable_variable_209_to_check)
);

// 变量节点210
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_210(
.clk(clk),
.rst(rst),
.initial_value(initial_value[210]),
.initial_value_enable(initial_value_enable[210]),
.initial_down(initial_down[210]),
.check_value_input(value_check_to_variable_210),
.check_enable_input(enable_check_to_variable_210),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_210_to_decision),
.value_variable_to_check(value_variable_210_to_check),
.variable_enable(enable_variable_210_to_check)
);

// 变量节点211
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_211(
.clk(clk),
.rst(rst),
.initial_value(initial_value[211]),
.initial_value_enable(initial_value_enable[211]),
.initial_down(initial_down[211]),
.check_value_input(value_check_to_variable_211),
.check_enable_input(enable_check_to_variable_211),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_211_to_decision),
.value_variable_to_check(value_variable_211_to_check),
.variable_enable(enable_variable_211_to_check)
);

// 变量节点212
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_212(
.clk(clk),
.rst(rst),
.initial_value(initial_value[212]),
.initial_value_enable(initial_value_enable[212]),
.initial_down(initial_down[212]),
.check_value_input(value_check_to_variable_212),
.check_enable_input(enable_check_to_variable_212),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_212_to_decision),
.value_variable_to_check(value_variable_212_to_check),
.variable_enable(enable_variable_212_to_check)
);

// 变量节点213
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_213(
.clk(clk),
.rst(rst),
.initial_value(initial_value[213]),
.initial_value_enable(initial_value_enable[213]),
.initial_down(initial_down[213]),
.check_value_input(value_check_to_variable_213),
.check_enable_input(enable_check_to_variable_213),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_213_to_decision),
.value_variable_to_check(value_variable_213_to_check),
.variable_enable(enable_variable_213_to_check)
);

// 变量节点214
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_214(
.clk(clk),
.rst(rst),
.initial_value(initial_value[214]),
.initial_value_enable(initial_value_enable[214]),
.initial_down(initial_down[214]),
.check_value_input(value_check_to_variable_214),
.check_enable_input(enable_check_to_variable_214),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_214_to_decision),
.value_variable_to_check(value_variable_214_to_check),
.variable_enable(enable_variable_214_to_check)
);

// 变量节点215
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_215(
.clk(clk),
.rst(rst),
.initial_value(initial_value[215]),
.initial_value_enable(initial_value_enable[215]),
.initial_down(initial_down[215]),
.check_value_input(value_check_to_variable_215),
.check_enable_input(enable_check_to_variable_215),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_215_to_decision),
.value_variable_to_check(value_variable_215_to_check),
.variable_enable(enable_variable_215_to_check)
);

// 变量节点216
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_216(
.clk(clk),
.rst(rst),
.initial_value(initial_value[216]),
.initial_value_enable(initial_value_enable[216]),
.initial_down(initial_down[216]),
.check_value_input(value_check_to_variable_216),
.check_enable_input(enable_check_to_variable_216),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_216_to_decision),
.value_variable_to_check(value_variable_216_to_check),
.variable_enable(enable_variable_216_to_check)
);

// 变量节点217
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_217(
.clk(clk),
.rst(rst),
.initial_value(initial_value[217]),
.initial_value_enable(initial_value_enable[217]),
.initial_down(initial_down[217]),
.check_value_input(value_check_to_variable_217),
.check_enable_input(enable_check_to_variable_217),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_217_to_decision),
.value_variable_to_check(value_variable_217_to_check),
.variable_enable(enable_variable_217_to_check)
);

// 变量节点218
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_218(
.clk(clk),
.rst(rst),
.initial_value(initial_value[218]),
.initial_value_enable(initial_value_enable[218]),
.initial_down(initial_down[218]),
.check_value_input(value_check_to_variable_218),
.check_enable_input(enable_check_to_variable_218),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_218_to_decision),
.value_variable_to_check(value_variable_218_to_check),
.variable_enable(enable_variable_218_to_check)
);

// 变量节点219
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_219(
.clk(clk),
.rst(rst),
.initial_value(initial_value[219]),
.initial_value_enable(initial_value_enable[219]),
.initial_down(initial_down[219]),
.check_value_input(value_check_to_variable_219),
.check_enable_input(enable_check_to_variable_219),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_219_to_decision),
.value_variable_to_check(value_variable_219_to_check),
.variable_enable(enable_variable_219_to_check)
);

// 变量节点220
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_220(
.clk(clk),
.rst(rst),
.initial_value(initial_value[220]),
.initial_value_enable(initial_value_enable[220]),
.initial_down(initial_down[220]),
.check_value_input(value_check_to_variable_220),
.check_enable_input(enable_check_to_variable_220),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_220_to_decision),
.value_variable_to_check(value_variable_220_to_check),
.variable_enable(enable_variable_220_to_check)
);

// 变量节点221
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_221(
.clk(clk),
.rst(rst),
.initial_value(initial_value[221]),
.initial_value_enable(initial_value_enable[221]),
.initial_down(initial_down[221]),
.check_value_input(value_check_to_variable_221),
.check_enable_input(enable_check_to_variable_221),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_221_to_decision),
.value_variable_to_check(value_variable_221_to_check),
.variable_enable(enable_variable_221_to_check)
);

// 变量节点222
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_222(
.clk(clk),
.rst(rst),
.initial_value(initial_value[222]),
.initial_value_enable(initial_value_enable[222]),
.initial_down(initial_down[222]),
.check_value_input(value_check_to_variable_222),
.check_enable_input(enable_check_to_variable_222),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_222_to_decision),
.value_variable_to_check(value_variable_222_to_check),
.variable_enable(enable_variable_222_to_check)
);

// 变量节点223
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_223(
.clk(clk),
.rst(rst),
.initial_value(initial_value[223]),
.initial_value_enable(initial_value_enable[223]),
.initial_down(initial_down[223]),
.check_value_input(value_check_to_variable_223),
.check_enable_input(enable_check_to_variable_223),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_223_to_decision),
.value_variable_to_check(value_variable_223_to_check),
.variable_enable(enable_variable_223_to_check)
);

// 变量节点224
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_224(
.clk(clk),
.rst(rst),
.initial_value(initial_value[224]),
.initial_value_enable(initial_value_enable[224]),
.initial_down(initial_down[224]),
.check_value_input(value_check_to_variable_224),
.check_enable_input(enable_check_to_variable_224),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_224_to_decision),
.value_variable_to_check(value_variable_224_to_check),
.variable_enable(enable_variable_224_to_check)
);

// 变量节点225
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_225(
.clk(clk),
.rst(rst),
.initial_value(initial_value[225]),
.initial_value_enable(initial_value_enable[225]),
.initial_down(initial_down[225]),
.check_value_input(value_check_to_variable_225),
.check_enable_input(enable_check_to_variable_225),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_225_to_decision),
.value_variable_to_check(value_variable_225_to_check),
.variable_enable(enable_variable_225_to_check)
);

// 变量节点226
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_226(
.clk(clk),
.rst(rst),
.initial_value(initial_value[226]),
.initial_value_enable(initial_value_enable[226]),
.initial_down(initial_down[226]),
.check_value_input(value_check_to_variable_226),
.check_enable_input(enable_check_to_variable_226),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_226_to_decision),
.value_variable_to_check(value_variable_226_to_check),
.variable_enable(enable_variable_226_to_check)
);

// 变量节点227
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_227(
.clk(clk),
.rst(rst),
.initial_value(initial_value[227]),
.initial_value_enable(initial_value_enable[227]),
.initial_down(initial_down[227]),
.check_value_input(value_check_to_variable_227),
.check_enable_input(enable_check_to_variable_227),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_227_to_decision),
.value_variable_to_check(value_variable_227_to_check),
.variable_enable(enable_variable_227_to_check)
);

// 变量节点228
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_228(
.clk(clk),
.rst(rst),
.initial_value(initial_value[228]),
.initial_value_enable(initial_value_enable[228]),
.initial_down(initial_down[228]),
.check_value_input(value_check_to_variable_228),
.check_enable_input(enable_check_to_variable_228),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_228_to_decision),
.value_variable_to_check(value_variable_228_to_check),
.variable_enable(enable_variable_228_to_check)
);

// 变量节点229
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_229(
.clk(clk),
.rst(rst),
.initial_value(initial_value[229]),
.initial_value_enable(initial_value_enable[229]),
.initial_down(initial_down[229]),
.check_value_input(value_check_to_variable_229),
.check_enable_input(enable_check_to_variable_229),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_229_to_decision),
.value_variable_to_check(value_variable_229_to_check),
.variable_enable(enable_variable_229_to_check)
);

// 变量节点230
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_230(
.clk(clk),
.rst(rst),
.initial_value(initial_value[230]),
.initial_value_enable(initial_value_enable[230]),
.initial_down(initial_down[230]),
.check_value_input(value_check_to_variable_230),
.check_enable_input(enable_check_to_variable_230),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_230_to_decision),
.value_variable_to_check(value_variable_230_to_check),
.variable_enable(enable_variable_230_to_check)
);

// 变量节点231
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_231(
.clk(clk),
.rst(rst),
.initial_value(initial_value[231]),
.initial_value_enable(initial_value_enable[231]),
.initial_down(initial_down[231]),
.check_value_input(value_check_to_variable_231),
.check_enable_input(enable_check_to_variable_231),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_231_to_decision),
.value_variable_to_check(value_variable_231_to_check),
.variable_enable(enable_variable_231_to_check)
);

// 变量节点232
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_232(
.clk(clk),
.rst(rst),
.initial_value(initial_value[232]),
.initial_value_enable(initial_value_enable[232]),
.initial_down(initial_down[232]),
.check_value_input(value_check_to_variable_232),
.check_enable_input(enable_check_to_variable_232),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_232_to_decision),
.value_variable_to_check(value_variable_232_to_check),
.variable_enable(enable_variable_232_to_check)
);

// 变量节点233
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_233(
.clk(clk),
.rst(rst),
.initial_value(initial_value[233]),
.initial_value_enable(initial_value_enable[233]),
.initial_down(initial_down[233]),
.check_value_input(value_check_to_variable_233),
.check_enable_input(enable_check_to_variable_233),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_233_to_decision),
.value_variable_to_check(value_variable_233_to_check),
.variable_enable(enable_variable_233_to_check)
);

// 变量节点234
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_234(
.clk(clk),
.rst(rst),
.initial_value(initial_value[234]),
.initial_value_enable(initial_value_enable[234]),
.initial_down(initial_down[234]),
.check_value_input(value_check_to_variable_234),
.check_enable_input(enable_check_to_variable_234),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_234_to_decision),
.value_variable_to_check(value_variable_234_to_check),
.variable_enable(enable_variable_234_to_check)
);

// 变量节点235
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_235(
.clk(clk),
.rst(rst),
.initial_value(initial_value[235]),
.initial_value_enable(initial_value_enable[235]),
.initial_down(initial_down[235]),
.check_value_input(value_check_to_variable_235),
.check_enable_input(enable_check_to_variable_235),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_235_to_decision),
.value_variable_to_check(value_variable_235_to_check),
.variable_enable(enable_variable_235_to_check)
);

// 变量节点236
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_236(
.clk(clk),
.rst(rst),
.initial_value(initial_value[236]),
.initial_value_enable(initial_value_enable[236]),
.initial_down(initial_down[236]),
.check_value_input(value_check_to_variable_236),
.check_enable_input(enable_check_to_variable_236),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_236_to_decision),
.value_variable_to_check(value_variable_236_to_check),
.variable_enable(enable_variable_236_to_check)
);

// 变量节点237
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_237(
.clk(clk),
.rst(rst),
.initial_value(initial_value[237]),
.initial_value_enable(initial_value_enable[237]),
.initial_down(initial_down[237]),
.check_value_input(value_check_to_variable_237),
.check_enable_input(enable_check_to_variable_237),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_237_to_decision),
.value_variable_to_check(value_variable_237_to_check),
.variable_enable(enable_variable_237_to_check)
);

// 变量节点238
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_238(
.clk(clk),
.rst(rst),
.initial_value(initial_value[238]),
.initial_value_enable(initial_value_enable[238]),
.initial_down(initial_down[238]),
.check_value_input(value_check_to_variable_238),
.check_enable_input(enable_check_to_variable_238),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_238_to_decision),
.value_variable_to_check(value_variable_238_to_check),
.variable_enable(enable_variable_238_to_check)
);

// 变量节点239
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_239(
.clk(clk),
.rst(rst),
.initial_value(initial_value[239]),
.initial_value_enable(initial_value_enable[239]),
.initial_down(initial_down[239]),
.check_value_input(value_check_to_variable_239),
.check_enable_input(enable_check_to_variable_239),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_239_to_decision),
.value_variable_to_check(value_variable_239_to_check),
.variable_enable(enable_variable_239_to_check)
);

// 变量节点240
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_240(
.clk(clk),
.rst(rst),
.initial_value(initial_value[240]),
.initial_value_enable(initial_value_enable[240]),
.initial_down(initial_down[240]),
.check_value_input(value_check_to_variable_240),
.check_enable_input(enable_check_to_variable_240),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_240_to_decision),
.value_variable_to_check(value_variable_240_to_check),
.variable_enable(enable_variable_240_to_check)
);

// 变量节点241
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_241(
.clk(clk),
.rst(rst),
.initial_value(initial_value[241]),
.initial_value_enable(initial_value_enable[241]),
.initial_down(initial_down[241]),
.check_value_input(value_check_to_variable_241),
.check_enable_input(enable_check_to_variable_241),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_241_to_decision),
.value_variable_to_check(value_variable_241_to_check),
.variable_enable(enable_variable_241_to_check)
);

// 变量节点242
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_242(
.clk(clk),
.rst(rst),
.initial_value(initial_value[242]),
.initial_value_enable(initial_value_enable[242]),
.initial_down(initial_down[242]),
.check_value_input(value_check_to_variable_242),
.check_enable_input(enable_check_to_variable_242),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_242_to_decision),
.value_variable_to_check(value_variable_242_to_check),
.variable_enable(enable_variable_242_to_check)
);

// 变量节点243
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_243(
.clk(clk),
.rst(rst),
.initial_value(initial_value[243]),
.initial_value_enable(initial_value_enable[243]),
.initial_down(initial_down[243]),
.check_value_input(value_check_to_variable_243),
.check_enable_input(enable_check_to_variable_243),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_243_to_decision),
.value_variable_to_check(value_variable_243_to_check),
.variable_enable(enable_variable_243_to_check)
);

// 变量节点244
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_244(
.clk(clk),
.rst(rst),
.initial_value(initial_value[244]),
.initial_value_enable(initial_value_enable[244]),
.initial_down(initial_down[244]),
.check_value_input(value_check_to_variable_244),
.check_enable_input(enable_check_to_variable_244),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_244_to_decision),
.value_variable_to_check(value_variable_244_to_check),
.variable_enable(enable_variable_244_to_check)
);

// 变量节点245
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_245(
.clk(clk),
.rst(rst),
.initial_value(initial_value[245]),
.initial_value_enable(initial_value_enable[245]),
.initial_down(initial_down[245]),
.check_value_input(value_check_to_variable_245),
.check_enable_input(enable_check_to_variable_245),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_245_to_decision),
.value_variable_to_check(value_variable_245_to_check),
.variable_enable(enable_variable_245_to_check)
);

// 变量节点246
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_246(
.clk(clk),
.rst(rst),
.initial_value(initial_value[246]),
.initial_value_enable(initial_value_enable[246]),
.initial_down(initial_down[246]),
.check_value_input(value_check_to_variable_246),
.check_enable_input(enable_check_to_variable_246),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_246_to_decision),
.value_variable_to_check(value_variable_246_to_check),
.variable_enable(enable_variable_246_to_check)
);

// 变量节点247
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_247(
.clk(clk),
.rst(rst),
.initial_value(initial_value[247]),
.initial_value_enable(initial_value_enable[247]),
.initial_down(initial_down[247]),
.check_value_input(value_check_to_variable_247),
.check_enable_input(enable_check_to_variable_247),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_247_to_decision),
.value_variable_to_check(value_variable_247_to_check),
.variable_enable(enable_variable_247_to_check)
);

// 变量节点248
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_248(
.clk(clk),
.rst(rst),
.initial_value(initial_value[248]),
.initial_value_enable(initial_value_enable[248]),
.initial_down(initial_down[248]),
.check_value_input(value_check_to_variable_248),
.check_enable_input(enable_check_to_variable_248),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_248_to_decision),
.value_variable_to_check(value_variable_248_to_check),
.variable_enable(enable_variable_248_to_check)
);

// 变量节点249
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_249(
.clk(clk),
.rst(rst),
.initial_value(initial_value[249]),
.initial_value_enable(initial_value_enable[249]),
.initial_down(initial_down[249]),
.check_value_input(value_check_to_variable_249),
.check_enable_input(enable_check_to_variable_249),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_249_to_decision),
.value_variable_to_check(value_variable_249_to_check),
.variable_enable(enable_variable_249_to_check)
);

// 变量节点250
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_250(
.clk(clk),
.rst(rst),
.initial_value(initial_value[250]),
.initial_value_enable(initial_value_enable[250]),
.initial_down(initial_down[250]),
.check_value_input(value_check_to_variable_250),
.check_enable_input(enable_check_to_variable_250),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_250_to_decision),
.value_variable_to_check(value_variable_250_to_check),
.variable_enable(enable_variable_250_to_check)
);

// 变量节点251
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_251(
.clk(clk),
.rst(rst),
.initial_value(initial_value[251]),
.initial_value_enable(initial_value_enable[251]),
.initial_down(initial_down[251]),
.check_value_input(value_check_to_variable_251),
.check_enable_input(enable_check_to_variable_251),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_251_to_decision),
.value_variable_to_check(value_variable_251_to_check),
.variable_enable(enable_variable_251_to_check)
);

// 变量节点252
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_252(
.clk(clk),
.rst(rst),
.initial_value(initial_value[252]),
.initial_value_enable(initial_value_enable[252]),
.initial_down(initial_down[252]),
.check_value_input(value_check_to_variable_252),
.check_enable_input(enable_check_to_variable_252),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_252_to_decision),
.value_variable_to_check(value_variable_252_to_check),
.variable_enable(enable_variable_252_to_check)
);

// 变量节点253
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_253(
.clk(clk),
.rst(rst),
.initial_value(initial_value[253]),
.initial_value_enable(initial_value_enable[253]),
.initial_down(initial_down[253]),
.check_value_input(value_check_to_variable_253),
.check_enable_input(enable_check_to_variable_253),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_253_to_decision),
.value_variable_to_check(value_variable_253_to_check),
.variable_enable(enable_variable_253_to_check)
);

// 变量节点254
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_254(
.clk(clk),
.rst(rst),
.initial_value(initial_value[254]),
.initial_value_enable(initial_value_enable[254]),
.initial_down(initial_down[254]),
.check_value_input(value_check_to_variable_254),
.check_enable_input(enable_check_to_variable_254),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_254_to_decision),
.value_variable_to_check(value_variable_254_to_check),
.variable_enable(enable_variable_254_to_check)
);

// 变量节点255
Variable_Node #(.weight(3), .length(6)) u_Variable_Node_255(
.clk(clk),
.rst(rst),
.initial_value(initial_value[255]),
.initial_value_enable(initial_value_enable[255]),
.initial_down(initial_down[255]),
.check_value_input(value_check_to_variable_255),
.check_enable_input(enable_check_to_variable_255),
.decision_down(decision_down),
.decoder_down(decoder_down),
.variable_value(value_variable_255_to_decision),
.value_variable_to_check(value_variable_255_to_check),
.variable_enable(enable_variable_255_to_check)
);



always@(*)begin
    // 调制结束，开始进行译码
    if(demodulation_down_to_decoder)begin
        prototype_sequence <= demodulation_prototype_sequence;
        initial_value_enable = 0-1;
    end
    else begin
        initial_value_enable = 0;
    end
    // 所有变量节点在初始化的时候信号是一致的，所以只需要对第一个变量节点进行讨论就行
    if(initial_down[0])begin
        demodulation_to_decoder_receive = 1;
    end
    else begin
        demodulation_to_decoder_receive = 0;
    end
end

// 校验部分与变量节点和校验节点的交互
always@(*)begin
    // 如果校验失败且迭代次数未到最大值,开始进行校验节点的更新
    if(decision_down & ~decision_success & ~decision_time_max) begin
        /*check_begin 可以是一位也可以是多位,看后面优化的时候怎么说*/
        check_begin = 1;
    end
    // 如果发现迭代次数到达最大值或者校验成功，那么译码结束
    if(decision_time_max || decision_success) begin
        /*这个也是,到底是一位还是多位优化时再考虑*/
        decoder_down = 1;
    end
    else decoder_down = 0;
end
// 将变量节点的enable值全部合并一下
assign decision_variable_enable[0] = enable_variable_0_to_check;
assign decision_variable_enable[1] = enable_variable_1_to_check;
assign decision_variable_enable[2] = enable_variable_2_to_check;
assign decision_variable_enable[3] = enable_variable_3_to_check;
assign decision_variable_enable[4] = enable_variable_4_to_check;
assign decision_variable_enable[5] = enable_variable_5_to_check;
assign decision_variable_enable[6] = enable_variable_6_to_check;
assign decision_variable_enable[7] = enable_variable_7_to_check;
assign decision_variable_enable[8] = enable_variable_8_to_check;
assign decision_variable_enable[9] = enable_variable_9_to_check;
assign decision_variable_enable[10] = enable_variable_10_to_check;
assign decision_variable_enable[11] = enable_variable_11_to_check;
assign decision_variable_enable[12] = enable_variable_12_to_check;
assign decision_variable_enable[13] = enable_variable_13_to_check;
assign decision_variable_enable[14] = enable_variable_14_to_check;
assign decision_variable_enable[15] = enable_variable_15_to_check;
assign decision_variable_enable[16] = enable_variable_16_to_check;
assign decision_variable_enable[17] = enable_variable_17_to_check;
assign decision_variable_enable[18] = enable_variable_18_to_check;
assign decision_variable_enable[19] = enable_variable_19_to_check;
assign decision_variable_enable[20] = enable_variable_20_to_check;
assign decision_variable_enable[21] = enable_variable_21_to_check;
assign decision_variable_enable[22] = enable_variable_22_to_check;
assign decision_variable_enable[23] = enable_variable_23_to_check;
assign decision_variable_enable[24] = enable_variable_24_to_check;
assign decision_variable_enable[25] = enable_variable_25_to_check;
assign decision_variable_enable[26] = enable_variable_26_to_check;
assign decision_variable_enable[27] = enable_variable_27_to_check;
assign decision_variable_enable[28] = enable_variable_28_to_check;
assign decision_variable_enable[29] = enable_variable_29_to_check;
assign decision_variable_enable[30] = enable_variable_30_to_check;
assign decision_variable_enable[31] = enable_variable_31_to_check;
assign decision_variable_enable[32] = enable_variable_32_to_check;
assign decision_variable_enable[33] = enable_variable_33_to_check;
assign decision_variable_enable[34] = enable_variable_34_to_check;
assign decision_variable_enable[35] = enable_variable_35_to_check;
assign decision_variable_enable[36] = enable_variable_36_to_check;
assign decision_variable_enable[37] = enable_variable_37_to_check;
assign decision_variable_enable[38] = enable_variable_38_to_check;
assign decision_variable_enable[39] = enable_variable_39_to_check;
assign decision_variable_enable[40] = enable_variable_40_to_check;
assign decision_variable_enable[41] = enable_variable_41_to_check;
assign decision_variable_enable[42] = enable_variable_42_to_check;
assign decision_variable_enable[43] = enable_variable_43_to_check;
assign decision_variable_enable[44] = enable_variable_44_to_check;
assign decision_variable_enable[45] = enable_variable_45_to_check;
assign decision_variable_enable[46] = enable_variable_46_to_check;
assign decision_variable_enable[47] = enable_variable_47_to_check;
assign decision_variable_enable[48] = enable_variable_48_to_check;
assign decision_variable_enable[49] = enable_variable_49_to_check;
assign decision_variable_enable[50] = enable_variable_50_to_check;
assign decision_variable_enable[51] = enable_variable_51_to_check;
assign decision_variable_enable[52] = enable_variable_52_to_check;
assign decision_variable_enable[53] = enable_variable_53_to_check;
assign decision_variable_enable[54] = enable_variable_54_to_check;
assign decision_variable_enable[55] = enable_variable_55_to_check;
assign decision_variable_enable[56] = enable_variable_56_to_check;
assign decision_variable_enable[57] = enable_variable_57_to_check;
assign decision_variable_enable[58] = enable_variable_58_to_check;
assign decision_variable_enable[59] = enable_variable_59_to_check;
assign decision_variable_enable[60] = enable_variable_60_to_check;
assign decision_variable_enable[61] = enable_variable_61_to_check;
assign decision_variable_enable[62] = enable_variable_62_to_check;
assign decision_variable_enable[63] = enable_variable_63_to_check;
assign decision_variable_enable[64] = enable_variable_64_to_check;
assign decision_variable_enable[65] = enable_variable_65_to_check;
assign decision_variable_enable[66] = enable_variable_66_to_check;
assign decision_variable_enable[67] = enable_variable_67_to_check;
assign decision_variable_enable[68] = enable_variable_68_to_check;
assign decision_variable_enable[69] = enable_variable_69_to_check;
assign decision_variable_enable[70] = enable_variable_70_to_check;
assign decision_variable_enable[71] = enable_variable_71_to_check;
assign decision_variable_enable[72] = enable_variable_72_to_check;
assign decision_variable_enable[73] = enable_variable_73_to_check;
assign decision_variable_enable[74] = enable_variable_74_to_check;
assign decision_variable_enable[75] = enable_variable_75_to_check;
assign decision_variable_enable[76] = enable_variable_76_to_check;
assign decision_variable_enable[77] = enable_variable_77_to_check;
assign decision_variable_enable[78] = enable_variable_78_to_check;
assign decision_variable_enable[79] = enable_variable_79_to_check;
assign decision_variable_enable[80] = enable_variable_80_to_check;
assign decision_variable_enable[81] = enable_variable_81_to_check;
assign decision_variable_enable[82] = enable_variable_82_to_check;
assign decision_variable_enable[83] = enable_variable_83_to_check;
assign decision_variable_enable[84] = enable_variable_84_to_check;
assign decision_variable_enable[85] = enable_variable_85_to_check;
assign decision_variable_enable[86] = enable_variable_86_to_check;
assign decision_variable_enable[87] = enable_variable_87_to_check;
assign decision_variable_enable[88] = enable_variable_88_to_check;
assign decision_variable_enable[89] = enable_variable_89_to_check;
assign decision_variable_enable[90] = enable_variable_90_to_check;
assign decision_variable_enable[91] = enable_variable_91_to_check;
assign decision_variable_enable[92] = enable_variable_92_to_check;
assign decision_variable_enable[93] = enable_variable_93_to_check;
assign decision_variable_enable[94] = enable_variable_94_to_check;
assign decision_variable_enable[95] = enable_variable_95_to_check;
assign decision_variable_enable[96] = enable_variable_96_to_check;
assign decision_variable_enable[97] = enable_variable_97_to_check;
assign decision_variable_enable[98] = enable_variable_98_to_check;
assign decision_variable_enable[99] = enable_variable_99_to_check;
assign decision_variable_enable[100] = enable_variable_100_to_check;
assign decision_variable_enable[101] = enable_variable_101_to_check;
assign decision_variable_enable[102] = enable_variable_102_to_check;
assign decision_variable_enable[103] = enable_variable_103_to_check;
assign decision_variable_enable[104] = enable_variable_104_to_check;
assign decision_variable_enable[105] = enable_variable_105_to_check;
assign decision_variable_enable[106] = enable_variable_106_to_check;
assign decision_variable_enable[107] = enable_variable_107_to_check;
assign decision_variable_enable[108] = enable_variable_108_to_check;
assign decision_variable_enable[109] = enable_variable_109_to_check;
assign decision_variable_enable[110] = enable_variable_110_to_check;
assign decision_variable_enable[111] = enable_variable_111_to_check;
assign decision_variable_enable[112] = enable_variable_112_to_check;
assign decision_variable_enable[113] = enable_variable_113_to_check;
assign decision_variable_enable[114] = enable_variable_114_to_check;
assign decision_variable_enable[115] = enable_variable_115_to_check;
assign decision_variable_enable[116] = enable_variable_116_to_check;
assign decision_variable_enable[117] = enable_variable_117_to_check;
assign decision_variable_enable[118] = enable_variable_118_to_check;
assign decision_variable_enable[119] = enable_variable_119_to_check;
assign decision_variable_enable[120] = enable_variable_120_to_check;
assign decision_variable_enable[121] = enable_variable_121_to_check;
assign decision_variable_enable[122] = enable_variable_122_to_check;
assign decision_variable_enable[123] = enable_variable_123_to_check;
assign decision_variable_enable[124] = enable_variable_124_to_check;
assign decision_variable_enable[125] = enable_variable_125_to_check;
assign decision_variable_enable[126] = enable_variable_126_to_check;
assign decision_variable_enable[127] = enable_variable_127_to_check;
assign decision_variable_enable[128] = enable_variable_128_to_check;
assign decision_variable_enable[129] = enable_variable_129_to_check;
assign decision_variable_enable[130] = enable_variable_130_to_check;
assign decision_variable_enable[131] = enable_variable_131_to_check;
assign decision_variable_enable[132] = enable_variable_132_to_check;
assign decision_variable_enable[133] = enable_variable_133_to_check;
assign decision_variable_enable[134] = enable_variable_134_to_check;
assign decision_variable_enable[135] = enable_variable_135_to_check;
assign decision_variable_enable[136] = enable_variable_136_to_check;
assign decision_variable_enable[137] = enable_variable_137_to_check;
assign decision_variable_enable[138] = enable_variable_138_to_check;
assign decision_variable_enable[139] = enable_variable_139_to_check;
assign decision_variable_enable[140] = enable_variable_140_to_check;
assign decision_variable_enable[141] = enable_variable_141_to_check;
assign decision_variable_enable[142] = enable_variable_142_to_check;
assign decision_variable_enable[143] = enable_variable_143_to_check;
assign decision_variable_enable[144] = enable_variable_144_to_check;
assign decision_variable_enable[145] = enable_variable_145_to_check;
assign decision_variable_enable[146] = enable_variable_146_to_check;
assign decision_variable_enable[147] = enable_variable_147_to_check;
assign decision_variable_enable[148] = enable_variable_148_to_check;
assign decision_variable_enable[149] = enable_variable_149_to_check;
assign decision_variable_enable[150] = enable_variable_150_to_check;
assign decision_variable_enable[151] = enable_variable_151_to_check;
assign decision_variable_enable[152] = enable_variable_152_to_check;
assign decision_variable_enable[153] = enable_variable_153_to_check;
assign decision_variable_enable[154] = enable_variable_154_to_check;
assign decision_variable_enable[155] = enable_variable_155_to_check;
assign decision_variable_enable[156] = enable_variable_156_to_check;
assign decision_variable_enable[157] = enable_variable_157_to_check;
assign decision_variable_enable[158] = enable_variable_158_to_check;
assign decision_variable_enable[159] = enable_variable_159_to_check;
assign decision_variable_enable[160] = enable_variable_160_to_check;
assign decision_variable_enable[161] = enable_variable_161_to_check;
assign decision_variable_enable[162] = enable_variable_162_to_check;
assign decision_variable_enable[163] = enable_variable_163_to_check;
assign decision_variable_enable[164] = enable_variable_164_to_check;
assign decision_variable_enable[165] = enable_variable_165_to_check;
assign decision_variable_enable[166] = enable_variable_166_to_check;
assign decision_variable_enable[167] = enable_variable_167_to_check;
assign decision_variable_enable[168] = enable_variable_168_to_check;
assign decision_variable_enable[169] = enable_variable_169_to_check;
assign decision_variable_enable[170] = enable_variable_170_to_check;
assign decision_variable_enable[171] = enable_variable_171_to_check;
assign decision_variable_enable[172] = enable_variable_172_to_check;
assign decision_variable_enable[173] = enable_variable_173_to_check;
assign decision_variable_enable[174] = enable_variable_174_to_check;
assign decision_variable_enable[175] = enable_variable_175_to_check;
assign decision_variable_enable[176] = enable_variable_176_to_check;
assign decision_variable_enable[177] = enable_variable_177_to_check;
assign decision_variable_enable[178] = enable_variable_178_to_check;
assign decision_variable_enable[179] = enable_variable_179_to_check;
assign decision_variable_enable[180] = enable_variable_180_to_check;
assign decision_variable_enable[181] = enable_variable_181_to_check;
assign decision_variable_enable[182] = enable_variable_182_to_check;
assign decision_variable_enable[183] = enable_variable_183_to_check;
assign decision_variable_enable[184] = enable_variable_184_to_check;
assign decision_variable_enable[185] = enable_variable_185_to_check;
assign decision_variable_enable[186] = enable_variable_186_to_check;
assign decision_variable_enable[187] = enable_variable_187_to_check;
assign decision_variable_enable[188] = enable_variable_188_to_check;
assign decision_variable_enable[189] = enable_variable_189_to_check;
assign decision_variable_enable[190] = enable_variable_190_to_check;
assign decision_variable_enable[191] = enable_variable_191_to_check;
assign decision_variable_enable[192] = enable_variable_192_to_check;
assign decision_variable_enable[193] = enable_variable_193_to_check;
assign decision_variable_enable[194] = enable_variable_194_to_check;
assign decision_variable_enable[195] = enable_variable_195_to_check;
assign decision_variable_enable[196] = enable_variable_196_to_check;
assign decision_variable_enable[197] = enable_variable_197_to_check;
assign decision_variable_enable[198] = enable_variable_198_to_check;
assign decision_variable_enable[199] = enable_variable_199_to_check;
assign decision_variable_enable[200] = enable_variable_200_to_check;
assign decision_variable_enable[201] = enable_variable_201_to_check;
assign decision_variable_enable[202] = enable_variable_202_to_check;
assign decision_variable_enable[203] = enable_variable_203_to_check;
assign decision_variable_enable[204] = enable_variable_204_to_check;
assign decision_variable_enable[205] = enable_variable_205_to_check;
assign decision_variable_enable[206] = enable_variable_206_to_check;
assign decision_variable_enable[207] = enable_variable_207_to_check;
assign decision_variable_enable[208] = enable_variable_208_to_check;
assign decision_variable_enable[209] = enable_variable_209_to_check;
assign decision_variable_enable[210] = enable_variable_210_to_check;
assign decision_variable_enable[211] = enable_variable_211_to_check;
assign decision_variable_enable[212] = enable_variable_212_to_check;
assign decision_variable_enable[213] = enable_variable_213_to_check;
assign decision_variable_enable[214] = enable_variable_214_to_check;
assign decision_variable_enable[215] = enable_variable_215_to_check;
assign decision_variable_enable[216] = enable_variable_216_to_check;
assign decision_variable_enable[217] = enable_variable_217_to_check;
assign decision_variable_enable[218] = enable_variable_218_to_check;
assign decision_variable_enable[219] = enable_variable_219_to_check;
assign decision_variable_enable[220] = enable_variable_220_to_check;
assign decision_variable_enable[221] = enable_variable_221_to_check;
assign decision_variable_enable[222] = enable_variable_222_to_check;
assign decision_variable_enable[223] = enable_variable_223_to_check;
assign decision_variable_enable[224] = enable_variable_224_to_check;
assign decision_variable_enable[225] = enable_variable_225_to_check;
assign decision_variable_enable[226] = enable_variable_226_to_check;
assign decision_variable_enable[227] = enable_variable_227_to_check;
assign decision_variable_enable[228] = enable_variable_228_to_check;
assign decision_variable_enable[229] = enable_variable_229_to_check;
assign decision_variable_enable[230] = enable_variable_230_to_check;
assign decision_variable_enable[231] = enable_variable_231_to_check;
assign decision_variable_enable[232] = enable_variable_232_to_check;
assign decision_variable_enable[233] = enable_variable_233_to_check;
assign decision_variable_enable[234] = enable_variable_234_to_check;
assign decision_variable_enable[235] = enable_variable_235_to_check;
assign decision_variable_enable[236] = enable_variable_236_to_check;
assign decision_variable_enable[237] = enable_variable_237_to_check;
assign decision_variable_enable[238] = enable_variable_238_to_check;
assign decision_variable_enable[239] = enable_variable_239_to_check;
assign decision_variable_enable[240] = enable_variable_240_to_check;
assign decision_variable_enable[241] = enable_variable_241_to_check;
assign decision_variable_enable[242] = enable_variable_242_to_check;
assign decision_variable_enable[243] = enable_variable_243_to_check;
assign decision_variable_enable[244] = enable_variable_244_to_check;
assign decision_variable_enable[245] = enable_variable_245_to_check;
assign decision_variable_enable[246] = enable_variable_246_to_check;
assign decision_variable_enable[247] = enable_variable_247_to_check;
assign decision_variable_enable[248] = enable_variable_248_to_check;
assign decision_variable_enable[249] = enable_variable_249_to_check;
assign decision_variable_enable[250] = enable_variable_250_to_check;
assign decision_variable_enable[251] = enable_variable_251_to_check;
assign decision_variable_enable[252] = enable_variable_252_to_check;
assign decision_variable_enable[253] = enable_variable_253_to_check;
assign decision_variable_enable[254] = enable_variable_254_to_check;
assign decision_variable_enable[255] = enable_variable_255_to_check;

integer i;
always@(posedge clk or negedge rst)begin
if(~rst)begin
i <= 0;
decision_state <= 0;
decision_down <= 0;
decision_success <= 0;
decision_information <= 0;
decision_times <= 0;
decision_result <= 0;
decision_time_max <= 0;
end
else begin
case(decision_state)
3'd0: begin
// 如果发现变量节点全部更新完毕,将变量节点的值进行判决然后计算
if(~decision_variable_enable == 0) begin
decision_information[0] <= value_variable_0_to_decision[5];
decision_information[1] <= value_variable_1_to_decision[5];
decision_information[2] <= value_variable_2_to_decision[5];
decision_information[3] <= value_variable_3_to_decision[5];
decision_information[4] <= value_variable_4_to_decision[5];
decision_information[5] <= value_variable_5_to_decision[5];
decision_information[6] <= value_variable_6_to_decision[5];
decision_information[7] <= value_variable_7_to_decision[5];
decision_information[8] <= value_variable_8_to_decision[5];
decision_information[9] <= value_variable_9_to_decision[5];
decision_information[10] <= value_variable_10_to_decision[5];
decision_information[11] <= value_variable_11_to_decision[5];
decision_information[12] <= value_variable_12_to_decision[5];
decision_information[13] <= value_variable_13_to_decision[5];
decision_information[14] <= value_variable_14_to_decision[5];
decision_information[15] <= value_variable_15_to_decision[5];
decision_information[16] <= value_variable_16_to_decision[5];
decision_information[17] <= value_variable_17_to_decision[5];
decision_information[18] <= value_variable_18_to_decision[5];
decision_information[19] <= value_variable_19_to_decision[5];
decision_information[20] <= value_variable_20_to_decision[5];
decision_information[21] <= value_variable_21_to_decision[5];
decision_information[22] <= value_variable_22_to_decision[5];
decision_information[23] <= value_variable_23_to_decision[5];
decision_information[24] <= value_variable_24_to_decision[5];
decision_information[25] <= value_variable_25_to_decision[5];
decision_information[26] <= value_variable_26_to_decision[5];
decision_information[27] <= value_variable_27_to_decision[5];
decision_information[28] <= value_variable_28_to_decision[5];
decision_information[29] <= value_variable_29_to_decision[5];
decision_information[30] <= value_variable_30_to_decision[5];
decision_information[31] <= value_variable_31_to_decision[5];
decision_information[32] <= value_variable_32_to_decision[5];
decision_information[33] <= value_variable_33_to_decision[5];
decision_information[34] <= value_variable_34_to_decision[5];
decision_information[35] <= value_variable_35_to_decision[5];
decision_information[36] <= value_variable_36_to_decision[5];
decision_information[37] <= value_variable_37_to_decision[5];
decision_information[38] <= value_variable_38_to_decision[5];
decision_information[39] <= value_variable_39_to_decision[5];
decision_information[40] <= value_variable_40_to_decision[5];
decision_information[41] <= value_variable_41_to_decision[5];
decision_information[42] <= value_variable_42_to_decision[5];
decision_information[43] <= value_variable_43_to_decision[5];
decision_information[44] <= value_variable_44_to_decision[5];
decision_information[45] <= value_variable_45_to_decision[5];
decision_information[46] <= value_variable_46_to_decision[5];
decision_information[47] <= value_variable_47_to_decision[5];
decision_information[48] <= value_variable_48_to_decision[5];
decision_information[49] <= value_variable_49_to_decision[5];
decision_information[50] <= value_variable_50_to_decision[5];
decision_information[51] <= value_variable_51_to_decision[5];
decision_information[52] <= value_variable_52_to_decision[5];
decision_information[53] <= value_variable_53_to_decision[5];
decision_information[54] <= value_variable_54_to_decision[5];
decision_information[55] <= value_variable_55_to_decision[5];
decision_information[56] <= value_variable_56_to_decision[5];
decision_information[57] <= value_variable_57_to_decision[5];
decision_information[58] <= value_variable_58_to_decision[5];
decision_information[59] <= value_variable_59_to_decision[5];
decision_information[60] <= value_variable_60_to_decision[5];
decision_information[61] <= value_variable_61_to_decision[5];
decision_information[62] <= value_variable_62_to_decision[5];
decision_information[63] <= value_variable_63_to_decision[5];
decision_information[64] <= value_variable_64_to_decision[5];
decision_information[65] <= value_variable_65_to_decision[5];
decision_information[66] <= value_variable_66_to_decision[5];
decision_information[67] <= value_variable_67_to_decision[5];
decision_information[68] <= value_variable_68_to_decision[5];
decision_information[69] <= value_variable_69_to_decision[5];
decision_information[70] <= value_variable_70_to_decision[5];
decision_information[71] <= value_variable_71_to_decision[5];
decision_information[72] <= value_variable_72_to_decision[5];
decision_information[73] <= value_variable_73_to_decision[5];
decision_information[74] <= value_variable_74_to_decision[5];
decision_information[75] <= value_variable_75_to_decision[5];
decision_information[76] <= value_variable_76_to_decision[5];
decision_information[77] <= value_variable_77_to_decision[5];
decision_information[78] <= value_variable_78_to_decision[5];
decision_information[79] <= value_variable_79_to_decision[5];
decision_information[80] <= value_variable_80_to_decision[5];
decision_information[81] <= value_variable_81_to_decision[5];
decision_information[82] <= value_variable_82_to_decision[5];
decision_information[83] <= value_variable_83_to_decision[5];
decision_information[84] <= value_variable_84_to_decision[5];
decision_information[85] <= value_variable_85_to_decision[5];
decision_information[86] <= value_variable_86_to_decision[5];
decision_information[87] <= value_variable_87_to_decision[5];
decision_information[88] <= value_variable_88_to_decision[5];
decision_information[89] <= value_variable_89_to_decision[5];
decision_information[90] <= value_variable_90_to_decision[5];
decision_information[91] <= value_variable_91_to_decision[5];
decision_information[92] <= value_variable_92_to_decision[5];
decision_information[93] <= value_variable_93_to_decision[5];
decision_information[94] <= value_variable_94_to_decision[5];
decision_information[95] <= value_variable_95_to_decision[5];
decision_information[96] <= value_variable_96_to_decision[5];
decision_information[97] <= value_variable_97_to_decision[5];
decision_information[98] <= value_variable_98_to_decision[5];
decision_information[99] <= value_variable_99_to_decision[5];
decision_information[100] <= value_variable_100_to_decision[5];
decision_information[101] <= value_variable_101_to_decision[5];
decision_information[102] <= value_variable_102_to_decision[5];
decision_information[103] <= value_variable_103_to_decision[5];
decision_information[104] <= value_variable_104_to_decision[5];
decision_information[105] <= value_variable_105_to_decision[5];
decision_information[106] <= value_variable_106_to_decision[5];
decision_information[107] <= value_variable_107_to_decision[5];
decision_information[108] <= value_variable_108_to_decision[5];
decision_information[109] <= value_variable_109_to_decision[5];
decision_information[110] <= value_variable_110_to_decision[5];
decision_information[111] <= value_variable_111_to_decision[5];
decision_information[112] <= value_variable_112_to_decision[5];
decision_information[113] <= value_variable_113_to_decision[5];
decision_information[114] <= value_variable_114_to_decision[5];
decision_information[115] <= value_variable_115_to_decision[5];
decision_information[116] <= value_variable_116_to_decision[5];
decision_information[117] <= value_variable_117_to_decision[5];
decision_information[118] <= value_variable_118_to_decision[5];
decision_information[119] <= value_variable_119_to_decision[5];
decision_information[120] <= value_variable_120_to_decision[5];
decision_information[121] <= value_variable_121_to_decision[5];
decision_information[122] <= value_variable_122_to_decision[5];
decision_information[123] <= value_variable_123_to_decision[5];
decision_information[124] <= value_variable_124_to_decision[5];
decision_information[125] <= value_variable_125_to_decision[5];
decision_information[126] <= value_variable_126_to_decision[5];
decision_information[127] <= value_variable_127_to_decision[5];
decision_information[128] <= value_variable_128_to_decision[5];
decision_information[129] <= value_variable_129_to_decision[5];
decision_information[130] <= value_variable_130_to_decision[5];
decision_information[131] <= value_variable_131_to_decision[5];
decision_information[132] <= value_variable_132_to_decision[5];
decision_information[133] <= value_variable_133_to_decision[5];
decision_information[134] <= value_variable_134_to_decision[5];
decision_information[135] <= value_variable_135_to_decision[5];
decision_information[136] <= value_variable_136_to_decision[5];
decision_information[137] <= value_variable_137_to_decision[5];
decision_information[138] <= value_variable_138_to_decision[5];
decision_information[139] <= value_variable_139_to_decision[5];
decision_information[140] <= value_variable_140_to_decision[5];
decision_information[141] <= value_variable_141_to_decision[5];
decision_information[142] <= value_variable_142_to_decision[5];
decision_information[143] <= value_variable_143_to_decision[5];
decision_information[144] <= value_variable_144_to_decision[5];
decision_information[145] <= value_variable_145_to_decision[5];
decision_information[146] <= value_variable_146_to_decision[5];
decision_information[147] <= value_variable_147_to_decision[5];
decision_information[148] <= value_variable_148_to_decision[5];
decision_information[149] <= value_variable_149_to_decision[5];
decision_information[150] <= value_variable_150_to_decision[5];
decision_information[151] <= value_variable_151_to_decision[5];
decision_information[152] <= value_variable_152_to_decision[5];
decision_information[153] <= value_variable_153_to_decision[5];
decision_information[154] <= value_variable_154_to_decision[5];
decision_information[155] <= value_variable_155_to_decision[5];
decision_information[156] <= value_variable_156_to_decision[5];
decision_information[157] <= value_variable_157_to_decision[5];
decision_information[158] <= value_variable_158_to_decision[5];
decision_information[159] <= value_variable_159_to_decision[5];
decision_information[160] <= value_variable_160_to_decision[5];
decision_information[161] <= value_variable_161_to_decision[5];
decision_information[162] <= value_variable_162_to_decision[5];
decision_information[163] <= value_variable_163_to_decision[5];
decision_information[164] <= value_variable_164_to_decision[5];
decision_information[165] <= value_variable_165_to_decision[5];
decision_information[166] <= value_variable_166_to_decision[5];
decision_information[167] <= value_variable_167_to_decision[5];
decision_information[168] <= value_variable_168_to_decision[5];
decision_information[169] <= value_variable_169_to_decision[5];
decision_information[170] <= value_variable_170_to_decision[5];
decision_information[171] <= value_variable_171_to_decision[5];
decision_information[172] <= value_variable_172_to_decision[5];
decision_information[173] <= value_variable_173_to_decision[5];
decision_information[174] <= value_variable_174_to_decision[5];
decision_information[175] <= value_variable_175_to_decision[5];
decision_information[176] <= value_variable_176_to_decision[5];
decision_information[177] <= value_variable_177_to_decision[5];
decision_information[178] <= value_variable_178_to_decision[5];
decision_information[179] <= value_variable_179_to_decision[5];
decision_information[180] <= value_variable_180_to_decision[5];
decision_information[181] <= value_variable_181_to_decision[5];
decision_information[182] <= value_variable_182_to_decision[5];
decision_information[183] <= value_variable_183_to_decision[5];
decision_information[184] <= value_variable_184_to_decision[5];
decision_information[185] <= value_variable_185_to_decision[5];
decision_information[186] <= value_variable_186_to_decision[5];
decision_information[187] <= value_variable_187_to_decision[5];
decision_information[188] <= value_variable_188_to_decision[5];
decision_information[189] <= value_variable_189_to_decision[5];
decision_information[190] <= value_variable_190_to_decision[5];
decision_information[191] <= value_variable_191_to_decision[5];
decision_information[192] <= value_variable_192_to_decision[5];
decision_information[193] <= value_variable_193_to_decision[5];
decision_information[194] <= value_variable_194_to_decision[5];
decision_information[195] <= value_variable_195_to_decision[5];
decision_information[196] <= value_variable_196_to_decision[5];
decision_information[197] <= value_variable_197_to_decision[5];
decision_information[198] <= value_variable_198_to_decision[5];
decision_information[199] <= value_variable_199_to_decision[5];
decision_information[200] <= value_variable_200_to_decision[5];
decision_information[201] <= value_variable_201_to_decision[5];
decision_information[202] <= value_variable_202_to_decision[5];
decision_information[203] <= value_variable_203_to_decision[5];
decision_information[204] <= value_variable_204_to_decision[5];
decision_information[205] <= value_variable_205_to_decision[5];
decision_information[206] <= value_variable_206_to_decision[5];
decision_information[207] <= value_variable_207_to_decision[5];
decision_information[208] <= value_variable_208_to_decision[5];
decision_information[209] <= value_variable_209_to_decision[5];
decision_information[210] <= value_variable_210_to_decision[5];
decision_information[211] <= value_variable_211_to_decision[5];
decision_information[212] <= value_variable_212_to_decision[5];
decision_information[213] <= value_variable_213_to_decision[5];
decision_information[214] <= value_variable_214_to_decision[5];
decision_information[215] <= value_variable_215_to_decision[5];
decision_information[216] <= value_variable_216_to_decision[5];
decision_information[217] <= value_variable_217_to_decision[5];
decision_information[218] <= value_variable_218_to_decision[5];
decision_information[219] <= value_variable_219_to_decision[5];
decision_information[220] <= value_variable_220_to_decision[5];
decision_information[221] <= value_variable_221_to_decision[5];
decision_information[222] <= value_variable_222_to_decision[5];
decision_information[223] <= value_variable_223_to_decision[5];
decision_information[224] <= value_variable_224_to_decision[5];
decision_information[225] <= value_variable_225_to_decision[5];
decision_information[226] <= value_variable_226_to_decision[5];
decision_information[227] <= value_variable_227_to_decision[5];
decision_information[228] <= value_variable_228_to_decision[5];
decision_information[229] <= value_variable_229_to_decision[5];
decision_information[230] <= value_variable_230_to_decision[5];
decision_information[231] <= value_variable_231_to_decision[5];
decision_information[232] <= value_variable_232_to_decision[5];
decision_information[233] <= value_variable_233_to_decision[5];
decision_information[234] <= value_variable_234_to_decision[5];
decision_information[235] <= value_variable_235_to_decision[5];
decision_information[236] <= value_variable_236_to_decision[5];
decision_information[237] <= value_variable_237_to_decision[5];
decision_information[238] <= value_variable_238_to_decision[5];
decision_information[239] <= value_variable_239_to_decision[5];
decision_information[240] <= value_variable_240_to_decision[5];
decision_information[241] <= value_variable_241_to_decision[5];
decision_information[242] <= value_variable_242_to_decision[5];
decision_information[243] <= value_variable_243_to_decision[5];
decision_information[244] <= value_variable_244_to_decision[5];
decision_information[245] <= value_variable_245_to_decision[5];
decision_information[246] <= value_variable_246_to_decision[5];
decision_information[247] <= value_variable_247_to_decision[5];
decision_information[248] <= value_variable_248_to_decision[5];
decision_information[249] <= value_variable_249_to_decision[5];
decision_information[250] <= value_variable_250_to_decision[5];
decision_information[251] <= value_variable_251_to_decision[5];
decision_information[252] <= value_variable_252_to_decision[5];
decision_information[253] <= value_variable_253_to_decision[5];
decision_information[254] <= value_variable_254_to_decision[5];
decision_information[255] <= value_variable_255_to_decision[5];
// 变更状态，开始进行校验
decision_state <= 3'd1;
end
end

// 开始校验
3'd1: begin
    // 一个周期完成校验
decision_result[0] <= decision_information[0] ^ decision_information[43] ^ decision_information[86] ^ decision_information[131] ^ decision_information[170] ^ decision_information[214];
decision_result[1] <= decision_information[1] ^ decision_information[42] ^ decision_information[87] ^ decision_information[132] ^ decision_information[173] ^ decision_information[215];
decision_result[2] <= decision_information[2] ^ decision_information[44] ^ decision_information[88] ^ decision_information[133] ^ decision_information[174] ^ decision_information[216];
decision_result[3] <= decision_information[3] ^ decision_information[45] ^ decision_information[89] ^ decision_information[134] ^ decision_information[175] ^ decision_information[217];
decision_result[4] <= decision_information[4] ^ decision_information[46] ^ decision_information[90] ^ decision_information[128] ^ decision_information[176] ^ decision_information[218];
decision_result[5] <= decision_information[5] ^ decision_information[47] ^ decision_information[91] ^ decision_information[135] ^ decision_information[177] ^ decision_information[219];
decision_result[6] <= decision_information[1] ^ decision_information[48] ^ decision_information[92] ^ decision_information[131] ^ decision_information[178] ^ decision_information[220];
decision_result[7] <= decision_information[6] ^ decision_information[47] ^ decision_information[93] ^ decision_information[136] ^ decision_information[179] ^ decision_information[221];
decision_result[8] <= decision_information[7] ^ decision_information[49] ^ decision_information[94] ^ decision_information[137] ^ decision_information[180] ^ decision_information[222];
decision_result[9] <= decision_information[8] ^ decision_information[50] ^ decision_information[95] ^ decision_information[138] ^ decision_information[179] ^ decision_information[223];
decision_result[10] <= decision_information[9] ^ decision_information[51] ^ decision_information[96] ^ decision_information[139] ^ decision_information[181] ^ decision_information[222];
decision_result[11] <= decision_information[10] ^ decision_information[52] ^ decision_information[97] ^ decision_information[140] ^ decision_information[182] ^ decision_information[224];
decision_result[12] <= decision_information[11] ^ decision_information[53] ^ decision_information[98] ^ decision_information[112] ^ decision_information[183] ^ decision_information[225];
decision_result[13] <= decision_information[12] ^ decision_information[54] ^ decision_information[99] ^ decision_information[141] ^ decision_information[184] ^ decision_information[226];
decision_result[14] <= decision_information[9] ^ decision_information[55] ^ decision_information[100] ^ decision_information[142] ^ decision_information[185] ^ decision_information[227];
decision_result[15] <= decision_information[12] ^ decision_information[56] ^ decision_information[101] ^ decision_information[143] ^ decision_information[186] ^ decision_information[217];
decision_result[16] <= decision_information[13] ^ decision_information[57] ^ decision_information[102] ^ decision_information[144] ^ decision_information[184] ^ decision_information[216];
decision_result[17] <= decision_information[14] ^ decision_information[58] ^ decision_information[102] ^ decision_information[145] ^ decision_information[187] ^ decision_information[228];
decision_result[18] <= decision_information[15] ^ decision_information[59] ^ decision_information[101] ^ decision_information[145] ^ decision_information[188] ^ decision_information[229];
decision_result[19] <= decision_information[16] ^ decision_information[60] ^ decision_information[92] ^ decision_information[146] ^ decision_information[186] ^ decision_information[230];
decision_result[20] <= decision_information[17] ^ decision_information[46] ^ decision_information[103] ^ decision_information[147] ^ decision_information[165] ^ decision_information[231];
decision_result[21] <= decision_information[18] ^ decision_information[61] ^ decision_information[104] ^ decision_information[132] ^ decision_information[188] ^ decision_information[218];
decision_result[22] <= decision_information[18] ^ decision_information[62] ^ decision_information[96] ^ decision_information[148] ^ decision_information[189] ^ decision_information[226];
decision_result[23] <= decision_information[19] ^ decision_information[55] ^ decision_information[94] ^ decision_information[149] ^ decision_information[190] ^ decision_information[232];
decision_result[24] <= decision_information[20] ^ decision_information[61] ^ decision_information[105] ^ decision_information[150] ^ decision_information[182] ^ decision_information[233];
decision_result[25] <= decision_information[21] ^ decision_information[50] ^ decision_information[106] ^ decision_information[137] ^ decision_information[191] ^ decision_information[234];
decision_result[26] <= decision_information[22] ^ decision_information[63] ^ decision_information[95] ^ decision_information[151] ^ decision_information[192] ^ decision_information[235];
decision_result[27] <= decision_information[23] ^ decision_information[64] ^ decision_information[107] ^ decision_information[152] ^ decision_information[193] ^ decision_information[225];
decision_result[28] <= decision_information[24] ^ decision_information[65] ^ decision_information[89] ^ decision_information[153] ^ decision_information[194] ^ decision_information[236];
decision_result[29] <= decision_information[11] ^ decision_information[66] ^ decision_information[104] ^ decision_information[154] ^ decision_information[180] ^ decision_information[237];
decision_result[30] <= decision_information[25] ^ decision_information[57] ^ decision_information[108] ^ decision_information[155] ^ decision_information[195] ^ decision_information[220];
decision_result[31] <= decision_information[26] ^ decision_information[59] ^ decision_information[109] ^ decision_information[156] ^ decision_information[195] ^ decision_information[236];
decision_result[32] <= decision_information[27] ^ decision_information[67] ^ decision_information[110] ^ decision_information[157] ^ decision_information[196] ^ decision_information[214];
decision_result[33] <= decision_information[28] ^ decision_information[49] ^ decision_information[111] ^ decision_information[158] ^ decision_information[189] ^ decision_information[225];
decision_result[34] <= decision_information[17] ^ decision_information[52] ^ decision_information[112] ^ decision_information[135] ^ decision_information[181] ^ decision_information[229];
decision_result[35] <= decision_information[0] ^ decision_information[64] ^ decision_information[113] ^ decision_information[135] ^ decision_information[197] ^ decision_information[230];
decision_result[36] <= decision_information[20] ^ decision_information[68] ^ decision_information[89] ^ decision_information[138] ^ decision_information[198] ^ decision_information[238];
decision_result[37] <= decision_information[19] ^ decision_information[67] ^ decision_information[101] ^ decision_information[129] ^ decision_information[189] ^ decision_information[213];
decision_result[38] <= decision_information[27] ^ decision_information[69] ^ decision_information[114] ^ decision_information[155] ^ decision_information[172] ^ decision_information[221];
decision_result[39] <= decision_information[21] ^ decision_information[70] ^ decision_information[115] ^ decision_information[146] ^ decision_information[199] ^ decision_information[239];
decision_result[40] <= decision_information[15] ^ decision_information[71] ^ decision_information[116] ^ decision_information[139] ^ decision_information[200] ^ decision_information[240];
decision_result[41] <= decision_information[20] ^ decision_information[64] ^ decision_information[90] ^ decision_information[142] ^ decision_information[201] ^ decision_information[241];
decision_result[42] <= decision_information[28] ^ decision_information[72] ^ decision_information[92] ^ decision_information[144] ^ decision_information[202] ^ decision_information[232];
decision_result[43] <= decision_information[29] ^ decision_information[73] ^ decision_information[117] ^ decision_information[143] ^ decision_information[176] ^ decision_information[219];
decision_result[44] <= decision_information[2] ^ decision_information[66] ^ decision_information[106] ^ decision_information[157] ^ decision_information[203] ^ decision_information[231];
decision_result[45] <= decision_information[30] ^ decision_information[62] ^ decision_information[118] ^ decision_information[159] ^ decision_information[195] ^ decision_information[227];
decision_result[46] <= decision_information[5] ^ decision_information[56] ^ decision_information[87] ^ decision_information[153] ^ decision_information[204] ^ decision_information[242];
decision_result[47] <= decision_information[31] ^ decision_information[51] ^ decision_information[119] ^ decision_information[143] ^ decision_information[198] ^ decision_information[228];
decision_result[48] <= decision_information[21] ^ decision_information[46] ^ decision_information[87] ^ decision_information[160] ^ decision_information[185] ^ decision_information[243];
decision_result[49] <= decision_information[32] ^ decision_information[74] ^ decision_information[119] ^ decision_information[136] ^ decision_information[183] ^ decision_information[240];
decision_result[50] <= decision_information[32] ^ decision_information[43] ^ decision_information[104] ^ decision_information[141] ^ decision_information[167] ^ decision_information[235];
decision_result[51] <= decision_information[7] ^ decision_information[75] ^ decision_information[119] ^ decision_information[150] ^ decision_information[205] ^ decision_information[244];
decision_result[52] <= decision_information[32] ^ decision_information[58] ^ decision_information[120] ^ decision_information[161] ^ decision_information[182] ^ decision_information[231];
decision_result[53] <= decision_information[33] ^ decision_information[63] ^ decision_information[121] ^ decision_information[152] ^ decision_information[174] ^ decision_information[243];
decision_result[54] <= decision_information[31] ^ decision_information[45] ^ decision_information[106] ^ decision_information[162] ^ decision_information[193] ^ decision_information[233];
decision_result[55] <= decision_information[34] ^ decision_information[62] ^ decision_information[103] ^ decision_information[134] ^ decision_information[177] ^ decision_information[245];
decision_result[56] <= decision_information[18] ^ decision_information[60] ^ decision_information[117] ^ decision_information[163] ^ decision_information[206] ^ decision_information[224];
decision_result[57] <= decision_information[8] ^ decision_information[76] ^ decision_information[86] ^ decision_information[100] ^ decision_information[172] ^ decision_information[228];
decision_result[58] <= decision_information[35] ^ decision_information[73] ^ decision_information[109] ^ decision_information[138] ^ decision_information[204] ^ decision_information[246];
decision_result[59] <= decision_information[24] ^ decision_information[77] ^ decision_information[99] ^ decision_information[146] ^ decision_information[193] ^ decision_information[246];
decision_result[60] <= decision_information[36] ^ decision_information[60] ^ decision_information[122] ^ decision_information[149] ^ decision_information[173] ^ decision_information[247];
decision_result[61] <= decision_information[7] ^ decision_information[44] ^ decision_information[114] ^ decision_information[151] ^ decision_information[202] ^ decision_information[242];
decision_result[62] <= decision_information[23] ^ decision_information[57] ^ decision_information[94] ^ decision_information[132] ^ decision_information[175] ^ decision_information[248];
decision_result[63] <= decision_information[22] ^ decision_information[78] ^ decision_information[113] ^ decision_information[156] ^ decision_information[207] ^ decision_information[217];
decision_result[64] <= decision_information[37] ^ decision_information[79] ^ decision_information[111] ^ decision_information[127] ^ decision_information[164] ^ decision_information[239];
decision_result[65] <= decision_information[24] ^ decision_information[58] ^ decision_information[114] ^ decision_information[160] ^ decision_information[197] ^ decision_information[249];
decision_result[66] <= decision_information[22] ^ decision_information[80] ^ decision_information[123] ^ decision_information[130] ^ decision_information[199] ^ decision_information[248];
decision_result[67] <= decision_information[31] ^ decision_information[81] ^ decision_information[91] ^ decision_information[164] ^ decision_information[180] ^ decision_information[223];
decision_result[68] <= decision_information[38] ^ decision_information[78] ^ decision_information[88] ^ decision_information[160] ^ decision_information[208] ^ decision_information[250];
decision_result[69] <= decision_information[38] ^ decision_information[48] ^ decision_information[110] ^ decision_information[139] ^ decision_information[177] ^ decision_information[212];
decision_result[70] <= decision_information[39] ^ decision_information[53] ^ decision_information[124] ^ decision_information[150] ^ decision_information[197] ^ decision_information[251];
decision_result[71] <= decision_information[40] ^ decision_information[61] ^ decision_information[110] ^ decision_information[158] ^ decision_information[191] ^ decision_information[227];
decision_result[72] <= decision_information[15] ^ decision_information[44] ^ decision_information[86] ^ decision_information[165] ^ decision_information[206] ^ decision_information[252];
decision_result[73] <= decision_information[6] ^ decision_information[77] ^ decision_information[96] ^ decision_information[156] ^ decision_information[209] ^ decision_information[216];
decision_result[74] <= decision_information[3] ^ decision_information[48] ^ decision_information[125] ^ decision_information[130] ^ decision_information[188] ^ decision_information[249];
decision_result[75] <= decision_information[26] ^ decision_information[81] ^ decision_information[103] ^ decision_information[141] ^ decision_information[200] ^ decision_information[234];
decision_result[76] <= decision_information[14] ^ decision_information[63] ^ decision_information[105] ^ decision_information[131] ^ decision_information[194] ^ decision_information[253];
decision_result[77] <= decision_information[37] ^ decision_information[50] ^ decision_information[107] ^ decision_information[140] ^ decision_information[205] ^ decision_information[245];
decision_result[78] <= decision_information[33] ^ decision_information[49] ^ decision_information[97] ^ decision_information[109] ^ decision_information[186] ^ decision_information[218];
decision_result[79] <= decision_information[39] ^ decision_information[78] ^ decision_information[111] ^ decision_information[163] ^ decision_information[210] ^ decision_information[242];
decision_result[80] <= decision_information[35] ^ decision_information[43] ^ decision_information[122] ^ decision_information[155] ^ decision_information[201] ^ decision_information[254];
decision_result[81] <= decision_information[13] ^ decision_information[76] ^ decision_information[124] ^ decision_information[148] ^ decision_information[201] ^ decision_information[234];
decision_result[82] <= decision_information[41] ^ decision_information[82] ^ decision_information[125] ^ decision_information[164] ^ decision_information[176] ^ decision_information[252];
decision_result[83] <= decision_information[29] ^ decision_information[55] ^ decision_information[126] ^ decision_information[140] ^ decision_information[203] ^ decision_information[220];
decision_result[84] <= decision_information[28] ^ decision_information[68] ^ decision_information[116] ^ decision_information[159] ^ decision_information[209] ^ decision_information[243];
decision_result[85] <= decision_information[25] ^ decision_information[77] ^ decision_information[127] ^ decision_information[129] ^ decision_information[183] ^ decision_information[250];
decision_result[86] <= decision_information[35] ^ decision_information[47] ^ decision_information[128] ^ decision_information[166] ^ decision_information[210] ^ decision_information[232];
decision_result[87] <= decision_information[29] ^ decision_information[71] ^ decision_information[98] ^ decision_information[162] ^ decision_information[208] ^ decision_information[239];
decision_result[88] <= decision_information[3] ^ decision_information[52] ^ decision_information[129] ^ decision_information[167] ^ decision_information[174] ^ decision_information[247];
decision_result[89] <= decision_information[37] ^ decision_information[65] ^ decision_information[122] ^ decision_information[147] ^ decision_information[196] ^ decision_information[219];
decision_result[90] <= decision_information[14] ^ decision_information[82] ^ decision_information[112] ^ decision_information[137] ^ decision_information[207] ^ decision_information[246];
decision_result[91] <= decision_information[4] ^ decision_information[71] ^ decision_information[121] ^ decision_information[161] ^ decision_information[190] ^ decision_information[230];
decision_result[92] <= decision_information[40] ^ decision_information[70] ^ decision_information[108] ^ decision_information[133] ^ decision_information[207] ^ decision_information[226];
decision_result[93] <= decision_information[8] ^ decision_information[72] ^ decision_information[118] ^ decision_information[161] ^ decision_information[199] ^ decision_information[247];
decision_result[94] <= decision_information[9] ^ decision_information[79] ^ decision_information[120] ^ decision_information[133] ^ decision_information[192] ^ decision_information[244];
decision_result[95] <= decision_information[16] ^ decision_information[59] ^ decision_information[124] ^ decision_information[168] ^ decision_information[208] ^ decision_information[255];
decision_result[96] <= decision_information[13] ^ decision_information[45] ^ decision_information[128] ^ decision_information[151] ^ decision_information[178] ^ decision_information[250];
decision_result[97] <= decision_information[41] ^ decision_information[54] ^ decision_information[88] ^ decision_information[149] ^ decision_information[211] ^ decision_information[240];
decision_result[98] <= decision_information[34] ^ decision_information[67] ^ decision_information[95] ^ decision_information[169] ^ decision_information[173] ^ decision_information[233];
decision_result[99] <= decision_information[2] ^ decision_information[83] ^ decision_information[117] ^ decision_information[168] ^ decision_information[212] ^ decision_information[215];
decision_result[100] <= decision_information[0] ^ decision_information[84] ^ decision_information[115] ^ decision_information[166] ^ decision_information[203] ^ decision_information[223];
decision_result[101] <= decision_information[4] ^ decision_information[80] ^ decision_information[99] ^ decision_information[158] ^ decision_information[181] ^ decision_information[221];
decision_result[102] <= decision_information[41] ^ decision_information[68] ^ decision_information[115] ^ decision_information[148] ^ decision_information[196] ^ decision_information[229];
decision_result[103] <= decision_information[38] ^ decision_information[73] ^ decision_information[102] ^ decision_information[165] ^ decision_information[192] ^ decision_information[251];
decision_result[104] <= decision_information[17] ^ decision_information[83] ^ decision_information[123] ^ decision_information[144] ^ decision_information[205] ^ decision_information[237];
decision_result[105] <= decision_information[19] ^ decision_information[83] ^ decision_information[93] ^ decision_information[170] ^ decision_information[204] ^ decision_information[249];
decision_result[106] <= decision_information[1] ^ decision_information[75] ^ decision_information[127] ^ decision_information[166] ^ decision_information[200] ^ decision_information[254];
decision_result[107] <= decision_information[10] ^ decision_information[54] ^ decision_information[118] ^ decision_information[162] ^ decision_information[213] ^ decision_information[222];
decision_result[108] <= decision_information[40] ^ decision_information[81] ^ decision_information[126] ^ decision_information[169] ^ decision_information[210] ^ decision_information[253];
decision_result[109] <= decision_information[34] ^ decision_information[85] ^ decision_information[116] ^ decision_information[154] ^ decision_information[184] ^ decision_information[236];
decision_result[110] <= decision_information[27] ^ decision_information[53] ^ decision_information[84] ^ decision_information[171] ^ decision_information[206] ^ decision_information[241];
decision_result[111] <= decision_information[10] ^ decision_information[74] ^ decision_information[108] ^ decision_information[153] ^ decision_information[187] ^ decision_information[255];
decision_result[112] <= decision_information[36] ^ decision_information[80] ^ decision_information[91] ^ decision_information[145] ^ decision_information[178] ^ decision_information[241];
decision_result[113] <= decision_information[26] ^ decision_information[69] ^ decision_information[107] ^ decision_information[163] ^ decision_information[213] ^ decision_information[238];
decision_result[114] <= decision_information[5] ^ decision_information[85] ^ decision_information[120] ^ decision_information[168] ^ decision_information[211] ^ decision_information[253];
decision_result[115] <= decision_information[42] ^ decision_information[69] ^ decision_information[123] ^ decision_information[159] ^ decision_information[194] ^ decision_information[251];
decision_result[116] <= decision_information[25] ^ decision_information[66] ^ decision_information[121] ^ decision_information[170] ^ decision_information[198] ^ decision_information[224];
decision_result[117] <= decision_information[11] ^ decision_information[56] ^ decision_information[130] ^ decision_information[142] ^ decision_information[179] ^ decision_information[214];
decision_result[118] <= decision_information[39] ^ decision_information[70] ^ decision_information[93] ^ decision_information[134] ^ decision_information[152] ^ decision_information[252];
decision_result[119] <= decision_information[12] ^ decision_information[79] ^ decision_information[105] ^ decision_information[172] ^ decision_information[190] ^ decision_information[215];
decision_result[120] <= decision_information[30] ^ decision_information[75] ^ decision_information[113] ^ decision_information[157] ^ decision_information[187] ^ decision_information[238];
decision_result[121] <= decision_information[16] ^ decision_information[74] ^ decision_information[90] ^ decision_information[169] ^ decision_information[209] ^ decision_information[237];
decision_result[122] <= decision_information[33] ^ decision_information[51] ^ decision_information[84] ^ decision_information[147] ^ decision_information[191] ^ decision_information[255];
decision_result[123] <= decision_information[42] ^ decision_information[82] ^ decision_information[100] ^ decision_information[136] ^ decision_information[202] ^ decision_information[245];
decision_result[124] <= decision_information[30] ^ decision_information[65] ^ decision_information[98] ^ decision_information[167] ^ decision_information[211] ^ decision_information[248];
decision_result[125] <= decision_information[6] ^ decision_information[72] ^ decision_information[126] ^ decision_information[171] ^ decision_information[212] ^ decision_information[235];
decision_result[126] <= decision_information[36] ^ decision_information[76] ^ decision_information[97] ^ decision_information[154] ^ decision_information[175] ^ decision_information[244];
decision_result[127] <= decision_information[23] ^ decision_information[85] ^ decision_information[125] ^ decision_information[171] ^ decision_information[185] ^ decision_information[254];

    decision_state <= 3'd2;
end

3'd2: begin
    // 校验成功
    if(decision_result == 0)begin
        decision_down <= 1;
        decision_success <= 1;
        // 让校验成功信号多保持一个周期
        decision_state <= 3'd4;
    end
    //此次校验没有成功
    else begin
        decision_down <= 1;
        decision_success <= 0;
        if(decision_times == 50) begin

            decision_time_max <= 1;
            decision_state <= 3'd4;
        end
        else begin 
            decision_times <= decision_times+1;
            decision_state <= 3'd3;
        end
    end
end

3'd3: begin
    decision_down <= 0;
    decision_time_max <= 0;
    decision_success <= 0;
    decision_state <= 3'd0;
end

// 拖延一周期时间
3'd4: begin
    decision_times <= 0;
    decision_state <= 3'd3;
end

endcase
end
end
endmodule
