/*
 * Author: neidong_fu
 * Time  : 2020/03/04
 * function: caculate ln(in0)
*/

module exp_log(
    // out = round(-2ln2*in * 2^8)
    input [6:0] in,         // in (1,6,0)
    output reg [14:0] out  // out(1,0,14)
    );
    
    always@(*) begin
        case(in)
            7'd   0:out =  15'd     0;
            7'd   1:out = -15'd   355;
            7'd   2:out = -15'd   710;
            7'd   3:out = -15'd  1065;
            7'd   4:out = -15'd  1420;
            7'd   5:out = -15'd  1774;
            7'd   6:out = -15'd  2129;
            7'd   7:out = -15'd  2484;
            7'd   8:out = -15'd  2839;
            7'd   9:out = -15'd  3194;
            7'd  10:out = -15'd  3549;
            7'd  11:out = -15'd  3904;
            7'd  12:out = -15'd  4259;
            7'd  13:out = -15'd  4614;
            7'd  14:out = -15'd  1968;
            7'd  15:out = -15'd  5323;
            7'd  16:out = -15'd  5678;
            7'd  17:out = -15'd  6033;
            7'd  18:out = -15'd  6388;
            7'd  19:out = -15'd  6743;
            7'd  20:out = -15'd  7098;
            7'd  21:out = -15'd  7453;
            7'd  22:out = -15'd  7808;
            7'd  23:out = -15'd  8163;
            7'd  24:out = -15'd  8517;
            7'd  25:out = -15'd  8872;
            7'd  26:out = -15'd  9227;
            7'd  27:out = -15'd  9582;
            7'd  28:out = -15'd  9937;
            7'd  29:out = -15'd 10292;
            7'd  30:out = -15'd 10647;
            7'd  31:out = -15'd 11002;
            7'd  32:out = -15'd 11357;
            7'd  33:out = -15'd 11711;
            7'd  34:out = -15'd 12066;
            7'd  35:out = -15'd 12421;
            7'd  36:out = -15'd 12776;
            7'd  37:out = -15'd 13131;
            7'd  38:out = -15'd 13486;
            7'd  39:out = -15'd 13841;
            7'd  40:out = -15'd 14196;
            7'd  41:out = -15'd 14551;
            7'd  42:out = -15'd 14905;
            7'd  43:out = -15'd 15260;
            7'd  44:out = -15'd 15615;
            7'd  45:out = -15'd 15970;
            7'd  46:out = -15'd 16325;
            7'd  47:out = -15'd 16384;
            7'd  48:out = -15'd 16384;
            7'd  49:out = -15'd 16384;
            7'd  50:out = -15'd 16384;
            7'd  51:out = -15'd 16384;
            7'd  52:out = -15'd 16384;
            7'd  53:out = -15'd 16384;
            7'd  54:out = -15'd 16384;
            7'd  55:out = -15'd 16384;
            7'd  56:out = -15'd 16384;
            7'd  57:out = -15'd 16384;
            7'd  58:out = -15'd 16384;
            7'd  59:out = -15'd 16384;
            7'd  60:out = -15'd 16384;
            7'd  61:out = -15'd 16384;
            7'd  62:out = -15'd 16384;
            7'd  63:out = -15'd 16384;
            7'd  64:out =  15'd 16383;        // index = 64(-64),1638. saturate to 16383
            7'd  65:out =  15'd 16383;
            7'd  66:out =  15'd 16383;
            7'd  67:out =  15'd 16383;
            7'd  68:out =  15'd 16383;
            7'd  69:out =  15'd 16383;
            7'd  70:out =  15'd 16383;
            7'd  71:out =  15'd 16383;
            7'd  72:out =  15'd 16383;
            7'd  73:out =  15'd 16383;
            7'd  74:out =  15'd 16383;
            7'd  75:out =  15'd 16383;
            7'd  76:out =  15'd 16383;
            7'd  77:out =  15'd 16383;
            7'd  78:out =  15'd 16383;
            7'd  79:out =  15'd 16383;
            7'd  80:out =  15'd 16383;
            7'd  81:out =  15'd 16383;
            7'd  82:out =  15'd 16325;
            7'd  83:out =  15'd 15970;
            7'd  84:out =  15'd 15615;
            7'd  85:out =  15'd 15260;
            7'd  86:out =  15'd 14905;
            7'd  87:out =  15'd 14551;
            7'd  88:out =  15'd 14196;
            7'd  89:out =  15'd 13841;
            7'd  90:out =  15'd 13486;
            7'd  91:out =  15'd 13131;
            7'd  92:out =  15'd 12776;
            7'd  93:out =  15'd 12421;
            7'd  94:out =  15'd 12066;
            7'd  95:out =  15'd 11711;
            7'd  96:out =  15'd 11357;
            7'd  97:out =  15'd 11002;
            7'd  98:out =  15'd 10647;
            7'd  99:out =  15'd 10292;
            7'd 100:out =  15'd 9937;
            7'd 101:out =  15'd 9582;
            7'd 102:out =  15'd 9227;
            7'd 103:out =  15'd 8872;
            7'd 104:out =  15'd 8517;
            7'd 105:out =  15'd 8163;
            7'd 106:out =  15'd 7808;
            7'd 107:out =  15'd 7453;
            7'd 108:out =  15'd 7098;
            7'd 109:out =  15'd 6743;
            7'd 110:out =  15'd 6388;
            7'd 111:out =  15'd 6033;
            7'd 112:out =  15'd 5678;
            7'd 113:out =  15'd 5323;
            7'd 114:out =  15'd 4968;
            7'd 115:out =  15'd 4614;
            7'd 116:out =  15'd 4259;
            7'd 117:out =  15'd 3904;
            7'd 118:out =  15'd 3549;
            7'd 119:out =  15'd 3194;
            7'd 120:out =  15'd 2839;
            7'd 121:out =  15'd 2484;
            7'd 122:out =  15'd 2129;
            7'd 123:out =  15'd 1774;
            7'd 124:out =  15'd 1420;
            7'd 125:out =  15'd 1065;
            7'd 126:out =  15'd 710;
            7'd 127:out =  15'd 355;           // index = 127(-1) ,355
            default: out = 15'd0;
        endcase
    end
    
endmodule
