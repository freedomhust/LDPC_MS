/*
 * Author: neidong_fu
 * Time  : 2020/03/04
 * function: caculate ln(mantissa)
*/

module man_log(
    // out = round(-2*ln(in/(2^10)) * 2^8)
    input [9:0] in,         // in (0,0,10)
    output reg [13:0] out  // out(0,0,14)
    );
    
    always@(*)begin
        case(in)
        10'd 1:out = 14'd 3549;
        10'd 2:out = 14'd 3194;
        10'd 3:out = 14'd 2986;
        10'd 4:out = 14'd 2839;
        10'd 5:out = 14'd 2725;
        10'd 6:out = 14'd 2632;
        10'd 7:out = 14'd 2553;
        10'd 8:out = 14'd 2484;
        10'd 9:out = 14'd 2424;
        10'd 10:out = 14'd 2370;
        10'd 11:out = 14'd 2321;
        10'd 12:out = 14'd 2277;
        10'd 13:out = 14'd 2236;
        10'd 14:out = 14'd 2198;
        10'd 15:out = 14'd 2162;
        10'd 16:out = 14'd 2129;
        10'd 17:out = 14'd 2098;
        10'd 18:out = 14'd 2069;
        10'd 19:out = 14'd 2041;
        10'd 20:out = 14'd 2015;
        10'd 21:out = 14'd 1990;
        10'd 22:out = 14'd 1966;
        10'd 23:out = 14'd 1944;
        10'd 24:out = 14'd 1922;
        10'd 25:out = 14'd 1901;
        10'd 26:out = 14'd 1881;
        10'd 27:out = 14'd 1861;
        10'd 28:out = 14'd 1843;
        10'd 29:out = 14'd 1825;
        10'd 30:out = 14'd 1808;
        10'd 31:out = 14'd 1791;
        10'd 32:out = 14'd 1774;
        10'd 33:out = 14'd 1759;
        10'd 34:out = 14'd 1743;
        10'd 35:out = 14'd 1729;
        10'd 36:out = 14'd 1714;
        10'd 37:out = 14'd 1700;
        10'd 38:out = 14'd 1686;
        10'd 39:out = 14'd 1673;
        10'd 40:out = 14'd 1660;
        10'd 41:out = 14'd 1648;
        10'd 42:out = 14'd 1635;
        10'd 43:out = 14'd 1623;
        10'd 44:out = 14'd 1611;
        10'd 45:out = 14'd 1600;
        10'd 46:out = 14'd 1589;
        10'd 47:out = 14'd 1578;
        10'd 48:out = 14'd 1567;
        10'd 49:out = 14'd 1556;
        10'd 50:out = 14'd 1546;
        10'd 51:out = 14'd 1536;
        10'd 52:out = 14'd 1526;
        10'd 53:out = 14'd 1516;
        10'd 54:out = 14'd 1507;
        10'd 55:out = 14'd 1497;
        10'd 56:out = 14'd 1488;
        10'd 57:out = 14'd 1479;
        10'd 58:out = 14'd 1470;
        10'd 59:out = 14'd 1461;
        10'd 60:out = 14'd 1453;
        10'd 61:out = 14'd 1444;
        10'd 62:out = 14'd 1436;
        10'd 63:out = 14'd 1428;
        10'd 64:out = 14'd 1420;
        10'd 65:out = 14'd 1412;
        10'd 66:out = 14'd 1404;
        10'd 67:out = 14'd 1396;
        10'd 68:out = 14'd 1389;
        10'd 69:out = 14'd 1381;
        10'd 70:out = 14'd 1374;
        10'd 71:out = 14'd 1366;
        10'd 72:out = 14'd 1359;
        10'd 73:out = 14'd 1352;
        10'd 74:out = 14'd 1345;
        10'd 75:out = 14'd 1338;
        10'd 76:out = 14'd 1332;
        10'd 77:out = 14'd 1325;
        10'd 78:out = 14'd 1318;
        10'd 79:out = 14'd 1312;
        10'd 80:out = 14'd 1305;
        10'd 81:out = 14'd 1299;
        10'd 82:out = 14'd 1293;
        10'd 83:out = 14'd 1286;
        10'd 84:out = 14'd 1280;
        10'd 85:out = 14'd 1274;
        10'd 86:out = 14'd 1268;
        10'd 87:out = 14'd 1262;
        10'd 88:out = 14'd 1257;
        10'd 89:out = 14'd 1251;
        10'd 90:out = 14'd 1245;
        10'd 91:out = 14'd 1239;
        10'd 92:out = 14'd 1234;
        10'd 93:out = 14'd 1228;
        10'd 94:out = 14'd 1223;
        10'd 95:out = 14'd 1217;
        10'd 96:out = 14'd 1212;
        10'd 97:out = 14'd 1207;
        10'd 98:out = 14'd 1201;
        10'd 99:out = 14'd 1196;
        10'd 100:out = 14'd 1191;
        10'd 101:out = 14'd 1186;
        10'd 102:out = 14'd 1181;
        10'd 103:out = 14'd 1176;
        10'd 104:out = 14'd 1171;
        10'd 105:out = 14'd 1166;
        10'd 106:out = 14'd 1161;
        10'd 107:out = 14'd 1156;
        10'd 108:out = 14'd 1152;
        10'd 109:out = 14'd 1147;
        10'd 110:out = 14'd 1142;
        10'd 111:out = 14'd 1138;
        10'd 112:out = 14'd 1133;
        10'd 113:out = 14'd 1128;
        10'd 114:out = 14'd 1124;
        10'd 115:out = 14'd 1120;
        10'd 116:out = 14'd 1115;
        10'd 117:out = 14'd 1111;
        10'd 118:out = 14'd 1106;
        10'd 119:out = 14'd 1102;
        10'd 120:out = 14'd 1098;
        10'd 121:out = 14'd 1093;
        10'd 122:out = 14'd 1089;
        10'd 123:out = 14'd 1085;
        10'd 124:out = 14'd 1081;
        10'd 125:out = 14'd 1077;
        10'd 126:out = 14'd 1073;
        10'd 127:out = 14'd 1069;
        10'd 128:out = 14'd 1065;
        10'd 129:out = 14'd 1061;
        10'd 130:out = 14'd 1057;
        10'd 131:out = 14'd 1053;
        10'd 132:out = 14'd 1049;
        10'd 133:out = 14'd 1045;
        10'd 134:out = 14'd 1041;
        10'd 135:out = 14'd 1037;
        10'd 136:out = 14'd 1034;
        10'd 137:out = 14'd 1030;
        10'd 138:out = 14'd 1026;
        10'd 139:out = 14'd 1022;
        10'd 140:out = 14'd 1019;
        10'd 141:out = 14'd 1015;
        10'd 142:out = 14'd 1012;
        10'd 143:out = 14'd 1008;
        10'd 144:out = 14'd 1004;
        10'd 145:out = 14'd 1001;
        10'd 146:out = 14'd 997;
        10'd 147:out = 14'd 994;
        10'd 148:out = 14'd 990;
        10'd 149:out = 14'd 987;
        10'd 150:out = 14'd 983;
        10'd 151:out = 14'd 980;
        10'd 152:out = 14'd 977;
        10'd 153:out = 14'd 973;
        10'd 154:out = 14'd 970;
        10'd 155:out = 14'd 967;
        10'd 156:out = 14'd 963;
        10'd 157:out = 14'd 960;
        10'd 158:out = 14'd 957;
        10'd 159:out = 14'd 954;
        10'd 160:out = 14'd 950;
        10'd 161:out = 14'd 947;
        10'd 162:out = 14'd 944;
        10'd 163:out = 14'd 941;
        10'd 164:out = 14'd 938;
        10'd 165:out = 14'd 935;
        10'd 166:out = 14'd 932;
        10'd 167:out = 14'd 929;
        10'd 168:out = 14'd 925;
        10'd 169:out = 14'd 922;
        10'd 170:out = 14'd 919;
        10'd 171:out = 14'd 916;
        10'd 172:out = 14'd 913;
        10'd 173:out = 14'd 910;
        10'd 174:out = 14'd 907;
        10'd 175:out = 14'd 905;
        10'd 176:out = 14'd 902;
        10'd 177:out = 14'd 899;
        10'd 178:out = 14'd 896;
        10'd 179:out = 14'd 893;
        10'd 180:out = 14'd 890;
        10'd 181:out = 14'd 887;
        10'd 182:out = 14'd 884;
        10'd 183:out = 14'd 882;
        10'd 184:out = 14'd 879;
        10'd 185:out = 14'd 876;
        10'd 186:out = 14'd 873;
        10'd 187:out = 14'd 871;
        10'd 188:out = 14'd 868;
        10'd 189:out = 14'd 865;
        10'd 190:out = 14'd 862;
        10'd 191:out = 14'd 860;
        10'd 192:out = 14'd 857;
        10'd 193:out = 14'd 854;
        10'd 194:out = 14'd 852;
        10'd 195:out = 14'd 849;
        10'd 196:out = 14'd 847;
        10'd 197:out = 14'd 844;
        10'd 198:out = 14'd 841;
        10'd 199:out = 14'd 839;
        10'd 200:out = 14'd 836;
        10'd 201:out = 14'd 834;
        10'd 202:out = 14'd 831;
        10'd 203:out = 14'd 829;
        10'd 204:out = 14'd 826;
        10'd 205:out = 14'd 824;
        10'd 206:out = 14'd 821;
        10'd 207:out = 14'd 819;
        10'd 208:out = 14'd 816;
        10'd 209:out = 14'd 814;
        10'd 210:out = 14'd 811;
        10'd 211:out = 14'd 809;
        10'd 212:out = 14'd 806;
        10'd 213:out = 14'd 804;
        10'd 214:out = 14'd 802;
        10'd 215:out = 14'd 799;
        10'd 216:out = 14'd 797;
        10'd 217:out = 14'd 794;
        10'd 218:out = 14'd 792;
        10'd 219:out = 14'd 790;
        10'd 220:out = 14'd 787;
        10'd 221:out = 14'd 785;
        10'd 222:out = 14'd 783;
        10'd 223:out = 14'd 780;
        10'd 224:out = 14'd 778;
        10'd 225:out = 14'd 776;
        10'd 226:out = 14'd 774;
        10'd 227:out = 14'd 771;
        10'd 228:out = 14'd 769;
        10'd 229:out = 14'd 767;
        10'd 230:out = 14'd 765;
        10'd 231:out = 14'd 762;
        10'd 232:out = 14'd 760;
        10'd 233:out = 14'd 758;
        10'd 234:out = 14'd 756;
        10'd 235:out = 14'd 754;
        10'd 236:out = 14'd 751;
        10'd 237:out = 14'd 749;
        10'd 238:out = 14'd 747;
        10'd 239:out = 14'd 745;
        10'd 240:out = 14'd 743;
        10'd 241:out = 14'd 741;
        10'd 242:out = 14'd 739;
        10'd 243:out = 14'd 736;
        10'd 244:out = 14'd 734;
        10'd 245:out = 14'd 732;
        10'd 246:out = 14'd 730;
        10'd 247:out = 14'd 728;
        10'd 248:out = 14'd 726;
        10'd 249:out = 14'd 724;
        10'd 250:out = 14'd 722;
        10'd 251:out = 14'd 720;
        10'd 252:out = 14'd 718;
        10'd 253:out = 14'd 716;
        10'd 254:out = 14'd 714;
        10'd 255:out = 14'd 712;
        10'd 256:out = 14'd 710;
        10'd 257:out = 14'd 708;
        10'd 258:out = 14'd 706;
        10'd 259:out = 14'd 704;
        10'd 260:out = 14'd 702;
        10'd 261:out = 14'd 700;
        10'd 262:out = 14'd 698;
        10'd 263:out = 14'd 696;
        10'd 264:out = 14'd 694;
        10'd 265:out = 14'd 692;
        10'd 266:out = 14'd 690;
        10'd 267:out = 14'd 688;
        10'd 268:out = 14'd 686;
        10'd 269:out = 14'd 684;
        10'd 270:out = 14'd 683;
        10'd 271:out = 14'd 681;
        10'd 272:out = 14'd 679;
        10'd 273:out = 14'd 677;
        10'd 274:out = 14'd 675;
        10'd 275:out = 14'd 673;
        10'd 276:out = 14'd 671;
        10'd 277:out = 14'd 669;
        10'd 278:out = 14'd 668;
        10'd 279:out = 14'd 666;
        10'd 280:out = 14'd 664;
        10'd 281:out = 14'd 662;
        10'd 282:out = 14'd 660;
        10'd 283:out = 14'd 658;
        10'd 284:out = 14'd 657;
        10'd 285:out = 14'd 655;
        10'd 286:out = 14'd 653;
        10'd 287:out = 14'd 651;
        10'd 288:out = 14'd 649;
        10'd 289:out = 14'd 648;
        10'd 290:out = 14'd 646;
        10'd 291:out = 14'd 644;
        10'd 292:out = 14'd 642;
        10'd 293:out = 14'd 641;
        10'd 294:out = 14'd 639;
        10'd 295:out = 14'd 637;
        10'd 296:out = 14'd 635;
        10'd 297:out = 14'd 634;
        10'd 298:out = 14'd 632;
        10'd 299:out = 14'd 630;
        10'd 300:out = 14'd 629;
        10'd 301:out = 14'd 627;
        10'd 302:out = 14'd 625;
        10'd 303:out = 14'd 623;
        10'd 304:out = 14'd 622;
        10'd 305:out = 14'd 620;
        10'd 306:out = 14'd 618;
        10'd 307:out = 14'd 617;
        10'd 308:out = 14'd 615;
        10'd 309:out = 14'd 613;
        10'd 310:out = 14'd 612;
        10'd 311:out = 14'd 610;
        10'd 312:out = 14'd 608;
        10'd 313:out = 14'd 607;
        10'd 314:out = 14'd 605;
        10'd 315:out = 14'd 604;
        10'd 316:out = 14'd 602;
        10'd 317:out = 14'd 600;
        10'd 318:out = 14'd 599;
        10'd 319:out = 14'd 597;
        10'd 320:out = 14'd 596;
        10'd 321:out = 14'd 594;
        10'd 322:out = 14'd 592;
        10'd 323:out = 14'd 591;
        10'd 324:out = 14'd 589;
        10'd 325:out = 14'd 588;
        10'd 326:out = 14'd 586;
        10'd 327:out = 14'd 584;
        10'd 328:out = 14'd 583;
        10'd 329:out = 14'd 581;
        10'd 330:out = 14'd 580;
        10'd 331:out = 14'd 578;
        10'd 332:out = 14'd 577;
        10'd 333:out = 14'd 575;
        10'd 334:out = 14'd 574;
        10'd 335:out = 14'd 572;
        10'd 336:out = 14'd 571;
        10'd 337:out = 14'd 569;
        10'd 338:out = 14'd 568;
        10'd 339:out = 14'd 566;
        10'd 340:out = 14'd 564;
        10'd 341:out = 14'd 563;
        10'd 342:out = 14'd 561;
        10'd 343:out = 14'd 560;
        10'd 344:out = 14'd 559;
        10'd 345:out = 14'd 557;
        10'd 346:out = 14'd 556;
        10'd 347:out = 14'd 554;
        10'd 348:out = 14'd 553;
        10'd 349:out = 14'd 551;
        10'd 350:out = 14'd 550;
        10'd 351:out = 14'd 548;
        10'd 352:out = 14'd 547;
        10'd 353:out = 14'd 545;
        10'd 354:out = 14'd 544;
        10'd 355:out = 14'd 542;
        10'd 356:out = 14'd 541;
        10'd 357:out = 14'd 540;
        10'd 358:out = 14'd 538;
        10'd 359:out = 14'd 537;
        10'd 360:out = 14'd 535;
        10'd 361:out = 14'd 534;
        10'd 362:out = 14'd 532;
        10'd 363:out = 14'd 531;
        10'd 364:out = 14'd 530;
        10'd 365:out = 14'd 528;
        10'd 366:out = 14'd 527;
        10'd 367:out = 14'd 525;
        10'd 368:out = 14'd 524;
        10'd 369:out = 14'd 523;
        10'd 370:out = 14'd 521;
        10'd 371:out = 14'd 520;
        10'd 372:out = 14'd 518;
        10'd 373:out = 14'd 517;
        10'd 374:out = 14'd 516;
        10'd 375:out = 14'd 514;
        10'd 376:out = 14'd 513;
        10'd 377:out = 14'd 512;
        10'd 378:out = 14'd 510;
        10'd 379:out = 14'd 509;
        10'd 380:out = 14'd 508;
        10'd 381:out = 14'd 506;
        10'd 382:out = 14'd 505;
        10'd 383:out = 14'd 504;
        10'd 384:out = 14'd 502;
        10'd 385:out = 14'd 501;
        10'd 386:out = 14'd 500;
        10'd 387:out = 14'd 498;
        10'd 388:out = 14'd 497;
        10'd 389:out = 14'd 496;
        10'd 390:out = 14'd 494;
        10'd 391:out = 14'd 493;
        10'd 392:out = 14'd 492;
        10'd 393:out = 14'd 490;
        10'd 394:out = 14'd 489;
        10'd 395:out = 14'd 488;
        10'd 396:out = 14'd 486;
        10'd 397:out = 14'd 485;
        10'd 398:out = 14'd 484;
        10'd 399:out = 14'd 483;
        10'd 400:out = 14'd 481;
        10'd 401:out = 14'd 480;
        10'd 402:out = 14'd 479;
        10'd 403:out = 14'd 477;
        10'd 404:out = 14'd 476;
        10'd 405:out = 14'd 475;
        10'd 406:out = 14'd 474;
        10'd 407:out = 14'd 472;
        10'd 408:out = 14'd 471;
        10'd 409:out = 14'd 470;
        10'd 410:out = 14'd 469;
        10'd 411:out = 14'd 467;
        10'd 412:out = 14'd 466;
        10'd 413:out = 14'd 465;
        10'd 414:out = 14'd 464;
        10'd 415:out = 14'd 462;
        10'd 416:out = 14'd 461;
        10'd 417:out = 14'd 460;
        10'd 418:out = 14'd 459;
        10'd 419:out = 14'd 458;
        10'd 420:out = 14'd 456;
        10'd 421:out = 14'd 455;
        10'd 422:out = 14'd 454;
        10'd 423:out = 14'd 453;
        10'd 424:out = 14'd 451;
        10'd 425:out = 14'd 450;
        10'd 426:out = 14'd 449;
        10'd 427:out = 14'd 448;
        10'd 428:out = 14'd 447;
        10'd 429:out = 14'd 445;
        10'd 430:out = 14'd 444;
        10'd 431:out = 14'd 443;
        10'd 432:out = 14'd 442;
        10'd 433:out = 14'd 441;
        10'd 434:out = 14'd 440;
        10'd 435:out = 14'd 438;
        10'd 436:out = 14'd 437;
        10'd 437:out = 14'd 436;
        10'd 438:out = 14'd 435;
        10'd 439:out = 14'd 434;
        10'd 440:out = 14'd 432;
        10'd 441:out = 14'd 431;
        10'd 442:out = 14'd 430;
        10'd 443:out = 14'd 429;
        10'd 444:out = 14'd 428;
        10'd 445:out = 14'd 427;
        10'd 446:out = 14'd 426;
        10'd 447:out = 14'd 424;
        10'd 448:out = 14'd 423;
        10'd 449:out = 14'd 422;
        10'd 450:out = 14'd 421;
        10'd 451:out = 14'd 420;
        10'd 452:out = 14'd 419;
        10'd 453:out = 14'd 418;
        10'd 454:out = 14'd 416;
        10'd 455:out = 14'd 415;
        10'd 456:out = 14'd 414;
        10'd 457:out = 14'd 413;
        10'd 458:out = 14'd 412;
        10'd 459:out = 14'd 411;
        10'd 460:out = 14'd 410;
        10'd 461:out = 14'd 409;
        10'd 462:out = 14'd 408;
        10'd 463:out = 14'd 406;
        10'd 464:out = 14'd 405;
        10'd 465:out = 14'd 404;
        10'd 466:out = 14'd 403;
        10'd 467:out = 14'd 402;
        10'd 468:out = 14'd 401;
        10'd 469:out = 14'd 400;
        10'd 470:out = 14'd 399;
        10'd 471:out = 14'd 398;
        10'd 472:out = 14'd 397;
        10'd 473:out = 14'd 395;
        10'd 474:out = 14'd 394;
        10'd 475:out = 14'd 393;
        10'd 476:out = 14'd 392;
        10'd 477:out = 14'd 391;
        10'd 478:out = 14'd 390;
        10'd 479:out = 14'd 389;
        10'd 480:out = 14'd 388;
        10'd 481:out = 14'd 387;
        10'd 482:out = 14'd 386;
        10'd 483:out = 14'd 385;
        10'd 484:out = 14'd 384;
        10'd 485:out = 14'd 383;
        10'd 486:out = 14'd 382;
        10'd 487:out = 14'd 381;
        10'd 488:out = 14'd 379;
        10'd 489:out = 14'd 378;
        10'd 490:out = 14'd 377;
        10'd 491:out = 14'd 376;
        10'd 492:out = 14'd 375;
        10'd 493:out = 14'd 374;
        10'd 494:out = 14'd 373;
        10'd 495:out = 14'd 372;
        10'd 496:out = 14'd 371;
        10'd 497:out = 14'd 370;
        10'd 498:out = 14'd 369;
        10'd 499:out = 14'd 368;
        10'd 500:out = 14'd 367;
        10'd 501:out = 14'd 366;
        10'd 502:out = 14'd 365;
        10'd 503:out = 14'd 364;
        10'd 504:out = 14'd 363;
        10'd 505:out = 14'd 362;
        10'd 506:out = 14'd 361;
        10'd 507:out = 14'd 360;
        10'd 508:out = 14'd 359;
        10'd 509:out = 14'd 358;
        10'd 510:out = 14'd 357;
        10'd 511:out = 14'd 356;
        10'd 512:out = 14'd 355;
        10'd 513:out = 14'd 354;
        10'd 514:out = 14'd 353;
        10'd 515:out = 14'd 352;
        10'd 516:out = 14'd 351;
        10'd 517:out = 14'd 350;
        10'd 518:out = 14'd 349;
        10'd 519:out = 14'd 348;
        10'd 520:out = 14'd 347;
        10'd 521:out = 14'd 346;
        10'd 522:out = 14'd 345;
        10'd 523:out = 14'd 344;
        10'd 524:out = 14'd 343;
        10'd 525:out = 14'd 342;
        10'd 526:out = 14'd 341;
        10'd 527:out = 14'd 340;
        10'd 528:out = 14'd 339;
        10'd 529:out = 14'd 338;
        10'd 530:out = 14'd 337;
        10'd 531:out = 14'd 336;
        10'd 532:out = 14'd 335;
        10'd 533:out = 14'd 334;
        10'd 534:out = 14'd 333;
        10'd 535:out = 14'd 332;
        10'd 536:out = 14'd 331;
        10'd 537:out = 14'd 330;
        10'd 538:out = 14'd 330;
        10'd 539:out = 14'd 329;
        10'd 540:out = 14'd 328;
        10'd 541:out = 14'd 327;
        10'd 542:out = 14'd 326;
        10'd 543:out = 14'd 325;
        10'd 544:out = 14'd 324;
        10'd 545:out = 14'd 323;
        10'd 546:out = 14'd 322;
        10'd 547:out = 14'd 321;
        10'd 548:out = 14'd 320;
        10'd 549:out = 14'd 319;
        10'd 550:out = 14'd 318;
        10'd 551:out = 14'd 317;
        10'd 552:out = 14'd 316;
        10'd 553:out = 14'd 315;
        10'd 554:out = 14'd 315;
        10'd 555:out = 14'd 314;
        10'd 556:out = 14'd 313;
        10'd 557:out = 14'd 312;
        10'd 558:out = 14'd 311;
        10'd 559:out = 14'd 310;
        10'd 560:out = 14'd 309;
        10'd 561:out = 14'd 308;
        10'd 562:out = 14'd 307;
        10'd 563:out = 14'd 306;
        10'd 564:out = 14'd 305;
        10'd 565:out = 14'd 304;
        10'd 566:out = 14'd 304;
        10'd 567:out = 14'd 303;
        10'd 568:out = 14'd 302;
        10'd 569:out = 14'd 301;
        10'd 570:out = 14'd 300;
        10'd 571:out = 14'd 299;
        10'd 572:out = 14'd 298;
        10'd 573:out = 14'd 297;
        10'd 574:out = 14'd 296;
        10'd 575:out = 14'd 295;
        10'd 576:out = 14'd 295;
        10'd 577:out = 14'd 294;
        10'd 578:out = 14'd 293;
        10'd 579:out = 14'd 292;
        10'd 580:out = 14'd 291;
        10'd 581:out = 14'd 290;
        10'd 582:out = 14'd 289;
        10'd 583:out = 14'd 288;
        10'd 584:out = 14'd 288;
        10'd 585:out = 14'd 287;
        10'd 586:out = 14'd 286;
        10'd 587:out = 14'd 285;
        10'd 588:out = 14'd 284;
        10'd 589:out = 14'd 283;
        10'd 590:out = 14'd 282;
        10'd 591:out = 14'd 281;
        10'd 592:out = 14'd 281;
        10'd 593:out = 14'd 280;
        10'd 594:out = 14'd 279;
        10'd 595:out = 14'd 278;
        10'd 596:out = 14'd 277;
        10'd 597:out = 14'd 276;
        10'd 598:out = 14'd 275;
        10'd 599:out = 14'd 275;
        10'd 600:out = 14'd 274;
        10'd 601:out = 14'd 273;
        10'd 602:out = 14'd 272;
        10'd 603:out = 14'd 271;
        10'd 604:out = 14'd 270;
        10'd 605:out = 14'd 269;
        10'd 606:out = 14'd 269;
        10'd 607:out = 14'd 268;
        10'd 608:out = 14'd 267;
        10'd 609:out = 14'd 266;
        10'd 610:out = 14'd 265;
        10'd 611:out = 14'd 264;
        10'd 612:out = 14'd 264;
        10'd 613:out = 14'd 263;
        10'd 614:out = 14'd 262;
        10'd 615:out = 14'd 261;
        10'd 616:out = 14'd 260;
        10'd 617:out = 14'd 259;
        10'd 618:out = 14'd 259;
        10'd 619:out = 14'd 258;
        10'd 620:out = 14'd 257;
        10'd 621:out = 14'd 256;
        10'd 622:out = 14'd 255;
        10'd 623:out = 14'd 254;
        10'd 624:out = 14'd 254;
        10'd 625:out = 14'd 253;
        10'd 626:out = 14'd 252;
        10'd 627:out = 14'd 251;
        10'd 628:out = 14'd 250;
        10'd 629:out = 14'd 250;
        10'd 630:out = 14'd 249;
        10'd 631:out = 14'd 248;
        10'd 632:out = 14'd 247;
        10'd 633:out = 14'd 246;
        10'd 634:out = 14'd 245;
        10'd 635:out = 14'd 245;
        10'd 636:out = 14'd 244;
        10'd 637:out = 14'd 243;
        10'd 638:out = 14'd 242;
        10'd 639:out = 14'd 241;
        10'd 640:out = 14'd 241;
        10'd 641:out = 14'd 240;
        10'd 642:out = 14'd 239;
        10'd 643:out = 14'd 238;
        10'd 644:out = 14'd 237;
        10'd 645:out = 14'd 237;
        10'd 646:out = 14'd 236;
        10'd 647:out = 14'd 235;
        10'd 648:out = 14'd 234;
        10'd 649:out = 14'd 233;
        10'd 650:out = 14'd 233;
        10'd 651:out = 14'd 232;
        10'd 652:out = 14'd 231;
        10'd 653:out = 14'd 230;
        10'd 654:out = 14'd 230;
        10'd 655:out = 14'd 229;
        10'd 656:out = 14'd 228;
        10'd 657:out = 14'd 227;
        10'd 658:out = 14'd 226;
        10'd 659:out = 14'd 226;
        10'd 660:out = 14'd 225;
        10'd 661:out = 14'd 224;
        10'd 662:out = 14'd 223;
        10'd 663:out = 14'd 223;
        10'd 664:out = 14'd 222;
        10'd 665:out = 14'd 221;
        10'd 666:out = 14'd 220;
        10'd 667:out = 14'd 219;
        10'd 668:out = 14'd 219;
        10'd 669:out = 14'd 218;
        10'd 670:out = 14'd 217;
        10'd 671:out = 14'd 216;
        10'd 672:out = 14'd 216;
        10'd 673:out = 14'd 215;
        10'd 674:out = 14'd 214;
        10'd 675:out = 14'd 213;
        10'd 676:out = 14'd 213;
        10'd 677:out = 14'd 212;
        10'd 678:out = 14'd 211;
        10'd 679:out = 14'd 210;
        10'd 680:out = 14'd 210;
        10'd 681:out = 14'd 209;
        10'd 682:out = 14'd 208;
        10'd 683:out = 14'd 207;
        10'd 684:out = 14'd 207;
        10'd 685:out = 14'd 206;
        10'd 686:out = 14'd 205;
        10'd 687:out = 14'd 204;
        10'd 688:out = 14'd 204;
        10'd 689:out = 14'd 203;
        10'd 690:out = 14'd 202;
        10'd 691:out = 14'd 201;
        10'd 692:out = 14'd 201;
        10'd 693:out = 14'd 200;
        10'd 694:out = 14'd 199;
        10'd 695:out = 14'd 198;
        10'd 696:out = 14'd 198;
        10'd 697:out = 14'd 197;
        10'd 698:out = 14'd 196;
        10'd 699:out = 14'd 195;
        10'd 700:out = 14'd 195;
        10'd 701:out = 14'd 194;
        10'd 702:out = 14'd 193;
        10'd 703:out = 14'd 193;
        10'd 704:out = 14'd 192;
        10'd 705:out = 14'd 191;
        10'd 706:out = 14'd 190;
        10'd 707:out = 14'd 190;
        10'd 708:out = 14'd 189;
        10'd 709:out = 14'd 188;
        10'd 710:out = 14'd 187;
        10'd 711:out = 14'd 187;
        10'd 712:out = 14'd 186;
        10'd 713:out = 14'd 185;
        10'd 714:out = 14'd 185;
        10'd 715:out = 14'd 184;
        10'd 716:out = 14'd 183;
        10'd 717:out = 14'd 182;
        10'd 718:out = 14'd 182;
        10'd 719:out = 14'd 181;
        10'd 720:out = 14'd 180;
        10'd 721:out = 14'd 180;
        10'd 722:out = 14'd 179;
        10'd 723:out = 14'd 178;
        10'd 724:out = 14'd 178;
        10'd 725:out = 14'd 177;
        10'd 726:out = 14'd 176;
        10'd 727:out = 14'd 175;
        10'd 728:out = 14'd 175;
        10'd 729:out = 14'd 174;
        10'd 730:out = 14'd 173;
        10'd 731:out = 14'd 173;
        10'd 732:out = 14'd 172;
        10'd 733:out = 14'd 171;
        10'd 734:out = 14'd 170;
        10'd 735:out = 14'd 170;
        10'd 736:out = 14'd 169;
        10'd 737:out = 14'd 168;
        10'd 738:out = 14'd 168;
        10'd 739:out = 14'd 167;
        10'd 740:out = 14'd 166;
        10'd 741:out = 14'd 166;
        10'd 742:out = 14'd 165;
        10'd 743:out = 14'd 164;
        10'd 744:out = 14'd 164;
        10'd 745:out = 14'd 163;
        10'd 746:out = 14'd 162;
        10'd 747:out = 14'd 161;
        10'd 748:out = 14'd 161;
        10'd 749:out = 14'd 160;
        10'd 750:out = 14'd 159;
        10'd 751:out = 14'd 159;
        10'd 752:out = 14'd 158;
        10'd 753:out = 14'd 157;
        10'd 754:out = 14'd 157;
        10'd 755:out = 14'd 156;
        10'd 756:out = 14'd 155;
        10'd 757:out = 14'd 155;
        10'd 758:out = 14'd 154;
        10'd 759:out = 14'd 153;
        10'd 760:out = 14'd 153;
        10'd 761:out = 14'd 152;
        10'd 762:out = 14'd 151;
        10'd 763:out = 14'd 151;
        10'd 764:out = 14'd 150;
        10'd 765:out = 14'd 149;
        10'd 766:out = 14'd 149;
        10'd 767:out = 14'd 148;
        10'd 768:out = 14'd 147;
        10'd 769:out = 14'd 147;
        10'd 770:out = 14'd 146;
        10'd 771:out = 14'd 145;
        10'd 772:out = 14'd 145;
        10'd 773:out = 14'd 144;
        10'd 774:out = 14'd 143;
        10'd 775:out = 14'd 143;
        10'd 776:out = 14'd 142;
        10'd 777:out = 14'd 141;
        10'd 778:out = 14'd 141;
        10'd 779:out = 14'd 140;
        10'd 780:out = 14'd 139;
        10'd 781:out = 14'd 139;
        10'd 782:out = 14'd 138;
        10'd 783:out = 14'd 137;
        10'd 784:out = 14'd 137;
        10'd 785:out = 14'd 136;
        10'd 786:out = 14'd 135;
        10'd 787:out = 14'd 135;
        10'd 788:out = 14'd 134;
        10'd 789:out = 14'd 133;
        10'd 790:out = 14'd 133;
        10'd 791:out = 14'd 132;
        10'd 792:out = 14'd 132;
        10'd 793:out = 14'd 131;
        10'd 794:out = 14'd 130;
        10'd 795:out = 14'd 130;
        10'd 796:out = 14'd 129;
        10'd 797:out = 14'd 128;
        10'd 798:out = 14'd 128;
        10'd 799:out = 14'd 127;
        10'd 800:out = 14'd 126;
        10'd 801:out = 14'd 126;
        10'd 802:out = 14'd 125;
        10'd 803:out = 14'd 124;
        10'd 804:out = 14'd 124;
        10'd 805:out = 14'd 123;
        10'd 806:out = 14'd 123;
        10'd 807:out = 14'd 122;
        10'd 808:out = 14'd 121;
        10'd 809:out = 14'd 121;
        10'd 810:out = 14'd 120;
        10'd 811:out = 14'd 119;
        10'd 812:out = 14'd 119;
        10'd 813:out = 14'd 118;
        10'd 814:out = 14'd 118;
        10'd 815:out = 14'd 117;
        10'd 816:out = 14'd 116;
        10'd 817:out = 14'd 116;
        10'd 818:out = 14'd 115;
        10'd 819:out = 14'd 114;
        10'd 820:out = 14'd 114;
        10'd 821:out = 14'd 113;
        10'd 822:out = 14'd 113;
        10'd 823:out = 14'd 112;
        10'd 824:out = 14'd 111;
        10'd 825:out = 14'd 111;
        10'd 826:out = 14'd 110;
        10'd 827:out = 14'd 109;
        10'd 828:out = 14'd 109;
        10'd 829:out = 14'd 108;
        10'd 830:out = 14'd 108;
        10'd 831:out = 14'd 107;
        10'd 832:out = 14'd 106;
        10'd 833:out = 14'd 106;
        10'd 834:out = 14'd 105;
        10'd 835:out = 14'd 104;
        10'd 836:out = 14'd 104;
        10'd 837:out = 14'd 103;
        10'd 838:out = 14'd 103;
        10'd 839:out = 14'd 102;
        10'd 840:out = 14'd 101;
        10'd 841:out = 14'd 101;
        10'd 842:out = 14'd 100;
        10'd 843:out = 14'd 100;
        10'd 844:out = 14'd 99;
        10'd 845:out = 14'd 98;
        10'd 846:out = 14'd 98;
        10'd 847:out = 14'd 97;
        10'd 848:out = 14'd 97;
        10'd 849:out = 14'd 96;
        10'd 850:out = 14'd 95;
        10'd 851:out = 14'd 95;
        10'd 852:out = 14'd 94;
        10'd 853:out = 14'd 94;
        10'd 854:out = 14'd 93;
        10'd 855:out = 14'd 92;
        10'd 856:out = 14'd 92;
        10'd 857:out = 14'd 91;
        10'd 858:out = 14'd 91;
        10'd 859:out = 14'd 90;
        10'd 860:out = 14'd 89;
        10'd 861:out = 14'd 89;
        10'd 862:out = 14'd 88;
        10'd 863:out = 14'd 88;
        10'd 864:out = 14'd 87;
        10'd 865:out = 14'd 86;
        10'd 866:out = 14'd 86;
        10'd 867:out = 14'd 85;
        10'd 868:out = 14'd 85;
        10'd 869:out = 14'd 84;
        10'd 870:out = 14'd 83;
        10'd 871:out = 14'd 83;
        10'd 872:out = 14'd 82;
        10'd 873:out = 14'd 82;
        10'd 874:out = 14'd 81;
        10'd 875:out = 14'd 81;
        10'd 876:out = 14'd 80;
        10'd 877:out = 14'd 79;
        10'd 878:out = 14'd 79;
        10'd 879:out = 14'd 78;
        10'd 880:out = 14'd 78;
        10'd 881:out = 14'd 77;
        10'd 882:out = 14'd 76;
        10'd 883:out = 14'd 76;
        10'd 884:out = 14'd 75;
        10'd 885:out = 14'd 75;
        10'd 886:out = 14'd 74;
        10'd 887:out = 14'd 74;
        10'd 888:out = 14'd 73;
        10'd 889:out = 14'd 72;
        10'd 890:out = 14'd 72;
        10'd 891:out = 14'd 71;
        10'd 892:out = 14'd 71;
        10'd 893:out = 14'd 70;
        10'd 894:out = 14'd 70;
        10'd 895:out = 14'd 69;
        10'd 896:out = 14'd 68;
        10'd 897:out = 14'd 68;
        10'd 898:out = 14'd 67;
        10'd 899:out = 14'd 67;
        10'd 900:out = 14'd 66;
        10'd 901:out = 14'd 66;
        10'd 902:out = 14'd 65;
        10'd 903:out = 14'd 64;
        10'd 904:out = 14'd 64;
        10'd 905:out = 14'd 63;
        10'd 906:out = 14'd 63;
        10'd 907:out = 14'd 62;
        10'd 908:out = 14'd 62;
        10'd 909:out = 14'd 61;
        10'd 910:out = 14'd 60;
        10'd 911:out = 14'd 60;
        10'd 912:out = 14'd 59;
        10'd 913:out = 14'd 59;
        10'd 914:out = 14'd 58;
        10'd 915:out = 14'd 58;
        10'd 916:out = 14'd 57;
        10'd 917:out = 14'd 57;
        10'd 918:out = 14'd 56;
        10'd 919:out = 14'd 55;
        10'd 920:out = 14'd 55;
        10'd 921:out = 14'd 54;
        10'd 922:out = 14'd 54;
        10'd 923:out = 14'd 53;
        10'd 924:out = 14'd 53;
        10'd 925:out = 14'd 52;
        10'd 926:out = 14'd 52;
        10'd 927:out = 14'd 51;
        10'd 928:out = 14'd 50;
        10'd 929:out = 14'd 50;
        10'd 930:out = 14'd 49;
        10'd 931:out = 14'd 49;
        10'd 932:out = 14'd 48;
        10'd 933:out = 14'd 48;
        10'd 934:out = 14'd 47;
        10'd 935:out = 14'd 47;
        10'd 936:out = 14'd 46;
        10'd 937:out = 14'd 45;
        10'd 938:out = 14'd 45;
        10'd 939:out = 14'd 44;
        10'd 940:out = 14'd 44;
        10'd 941:out = 14'd 43;
        10'd 942:out = 14'd 43;
        10'd 943:out = 14'd 42;
        10'd 944:out = 14'd 42;
        10'd 945:out = 14'd 41;
        10'd 946:out = 14'd 41;
        10'd 947:out = 14'd 40;
        10'd 948:out = 14'd 39;
        10'd 949:out = 14'd 39;
        10'd 950:out = 14'd 38;
        10'd 951:out = 14'd 38;
        10'd 952:out = 14'd 37;
        10'd 953:out = 14'd 37;
        10'd 954:out = 14'd 36;
        10'd 955:out = 14'd 36;
        10'd 956:out = 14'd 35;
        10'd 957:out = 14'd 35;
        10'd 958:out = 14'd 34;
        10'd 959:out = 14'd 34;
        10'd 960:out = 14'd 33;
        10'd 961:out = 14'd 33;
        10'd 962:out = 14'd 32;
        10'd 963:out = 14'd 31;
        10'd 964:out = 14'd 31;
        10'd 965:out = 14'd 30;
        10'd 966:out = 14'd 30;
        10'd 967:out = 14'd 29;
        10'd 968:out = 14'd 29;
        10'd 969:out = 14'd 28;
        10'd 970:out = 14'd 28;
        10'd 971:out = 14'd 27;
        10'd 972:out = 14'd 27;
        10'd 973:out = 14'd 26;
        10'd 974:out = 14'd 26;
        10'd 975:out = 14'd 25;
        10'd 976:out = 14'd 25;
        10'd 977:out = 14'd 24;
        10'd 978:out = 14'd 24;
        10'd 979:out = 14'd 23;
        10'd 980:out = 14'd 22;
        10'd 981:out = 14'd 22;
        10'd 982:out = 14'd 21;
        10'd 983:out = 14'd 21;
        10'd 984:out = 14'd 20;
        10'd 985:out = 14'd 20;
        10'd 986:out = 14'd 19;
        10'd 987:out = 14'd 19;
        10'd 988:out = 14'd 18;
        10'd 989:out = 14'd 18;
        10'd 990:out = 14'd 17;
        10'd 991:out = 14'd 17;
        10'd 992:out = 14'd 16;
        10'd 993:out = 14'd 16;
        10'd 994:out = 14'd 15;
        10'd 995:out = 14'd 15;
        10'd 996:out = 14'd 14;
        10'd 997:out = 14'd 14;
        10'd 998:out = 14'd 13;
        10'd 999:out = 14'd 13;
        10'd 1000:out = 14'd 12;
        10'd 1001:out = 14'd 12;
        10'd 1002:out = 14'd 11;
        10'd 1003:out = 14'd 11;
        10'd 1004:out = 14'd 10;
        10'd 1005:out = 14'd 10;
        10'd 1006:out = 14'd 9;
        10'd 1007:out = 14'd 9;
        10'd 1008:out = 14'd 8;
        10'd 1009:out = 14'd 8;
        10'd 1010:out = 14'd 7;
        10'd 1011:out = 14'd 7;
        10'd 1012:out = 14'd 6;
        10'd 1013:out = 14'd 6;
        10'd 1014:out = 14'd 5;
        10'd 1015:out = 14'd 5;
        10'd 1016:out = 14'd 4;
        10'd 1017:out = 14'd 4;
        10'd 1018:out = 14'd 3;
        10'd 1019:out = 14'd 3;
        10'd 1020:out = 14'd 2;
        10'd 1021:out = 14'd 2;
        10'd 1022:out = 14'd 1;
        10'd 1023:out = 14'd 1;
            default  :out = 14'd    0;
        endcase
    end
    
endmodule
